//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.09 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Sat Jan 28 18:45:28 2023

module Gowin_SP (dout, clk, oce, ce, reset, wre, ad, din);

output [15:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [14:0] ad;
input [15:0] din;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire [26:0] spx9_inst_0_dout_w;
wire [8:0] spx9_inst_0_dout;
wire [26:0] spx9_inst_1_dout_w;
wire [8:0] spx9_inst_1_dout;
wire [26:0] spx9_inst_2_dout_w;
wire [8:0] spx9_inst_2_dout;
wire [26:0] spx9_inst_3_dout_w;
wire [8:0] spx9_inst_3_dout;
wire [26:0] spx9_inst_4_dout_w;
wire [8:0] spx9_inst_4_dout;
wire [26:0] spx9_inst_5_dout_w;
wire [8:0] spx9_inst_5_dout;
wire [26:0] spx9_inst_6_dout_w;
wire [8:0] spx9_inst_6_dout;
wire [26:0] spx9_inst_7_dout_w;
wire [8:0] spx9_inst_7_dout;
wire [30:0] sp_inst_8_dout_w;
wire [9:9] sp_inst_8_dout;
wire [30:0] sp_inst_9_dout_w;
wire [10:10] sp_inst_9_dout;
wire [30:0] sp_inst_10_dout_w;
wire [11:11] sp_inst_10_dout;
wire [30:0] sp_inst_11_dout_w;
wire [12:12] sp_inst_11_dout;
wire [30:0] sp_inst_12_dout_w;
wire [13:13] sp_inst_12_dout;
wire [30:0] sp_inst_13_dout_w;
wire [14:14] sp_inst_13_dout;
wire [30:0] sp_inst_14_dout_w;
wire [15:15] sp_inst_14_dout;
wire [29:0] sp_inst_15_dout_w;
wire [1:0] sp_inst_15_dout;
wire [29:0] sp_inst_16_dout_w;
wire [3:2] sp_inst_16_dout;
wire [29:0] sp_inst_17_dout_w;
wire [5:4] sp_inst_17_dout;
wire [29:0] sp_inst_18_dout_w;
wire [7:6] sp_inst_18_dout;
wire [29:0] sp_inst_19_dout_w;
wire [9:8] sp_inst_19_dout;
wire [29:0] sp_inst_20_dout_w;
wire [11:10] sp_inst_20_dout;
wire [29:0] sp_inst_21_dout_w;
wire [13:12] sp_inst_21_dout;
wire [29:0] sp_inst_22_dout_w;
wire [15:14] sp_inst_22_dout;
wire [15:0] sp_inst_23_dout_w;
wire [15:0] sp_inst_23_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_16;
wire mux_o_17;
wire mux_o_20;
wire mux_o_21;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_39;
wire mux_o_40;
wire mux_o_43;
wire mux_o_44;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_62;
wire mux_o_63;
wire mux_o_66;
wire mux_o_67;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_85;
wire mux_o_86;
wire mux_o_89;
wire mux_o_90;
wire mux_o_102;
wire mux_o_103;
wire mux_o_104;
wire mux_o_105;
wire mux_o_108;
wire mux_o_109;
wire mux_o_112;
wire mux_o_113;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_131;
wire mux_o_132;
wire mux_o_135;
wire mux_o_136;
wire mux_o_148;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_154;
wire mux_o_155;
wire mux_o_158;
wire mux_o_159;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_177;
wire mux_o_178;
wire mux_o_181;
wire mux_o_182;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_200;
wire mux_o_201;
wire mux_o_204;
wire mux_o_205;
wire mux_o_217;
wire mux_o_229;
wire mux_o_241;
wire mux_o_253;
wire mux_o_265;
wire mux_o_277;
wire mux_o_289;
wire ce_w;
wire gw_vcc;
wire gw_gnd;

assign ce_w = ~wre & ce;
assign gw_vcc = 1'b1;
assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_1.INIT = 16'h0002;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_2.INIT = 16'h0004;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_3.INIT = 16'h0008;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_4.INIT = 16'h0010;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_5.INIT = 16'h0020;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_6.INIT = 16'h0040;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(ad[11]),
  .I1(ad[12]),
  .I2(ad[13]),
  .I3(ad[14])
);
defparam lut_inst_7.INIT = 16'h0080;
LUT5 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[10]),
  .I1(ad[11]),
  .I2(ad[12]),
  .I3(ad[13]),
  .I4(ad[14])
);
defparam lut_inst_8.INIT = 32'h01000000;
SPX9 spx9_inst_0 (
    .DO({spx9_inst_0_dout_w[26:0],spx9_inst_0_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_0}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_0.READ_MODE = 1'b0;
defparam spx9_inst_0.WRITE_MODE = 2'b00;
defparam spx9_inst_0.BIT_WIDTH = 9;
defparam spx9_inst_0.BLK_SEL = 3'b001;
defparam spx9_inst_0.RESET_MODE = "SYNC";
defparam spx9_inst_0.INIT_RAM_00 = 288'hEAD499C2BC441588A351A8CC44110904C46241A0D06A341A0D068341A0D0683412090462;
defparam spx9_inst_0.INIT_RAM_01 = 288'h6A24FE37087BBD9EAF479BCDED088DCF6BF60B0DCAE571B8DC6E370B85BEC160B8DC6E36;
defparam spx9_inst_0.INIT_RAM_02 = 288'hEAF57EDD5CA5D32995CAE572B95CADD2260FB642DD50BA66B41E7128EBD58CDD824E2914;
defparam spx9_inst_0.INIT_RAM_03 = 288'h6D36974995CB69B4DA4CA60F0997D46DF4B95CAE9B4DA4CA6532581B8DC2DF6EAF57EDD5;
defparam spx9_inst_0.INIT_RAM_04 = 288'h2C1E06FF6FB7D82E784C9E132B95CA6532B95D36972B96D26574FA6D36974992B960B078;
defparam spx9_inst_0.INIT_RAM_05 = 288'h482C5E51389C4E26F27944A6754BA6576BB5CA6D42C16FB757ABD5EAF57EBF6FB7D82C37;
defparam spx9_inst_0.INIT_RAM_06 = 288'h20988C48341A0D468341A0D068351A0D068341A0905B7DB656E9549A44E2733893456270;
defparam spx9_inst_0.INIT_RAM_07 = 288'hA96536BD5FB7D82E372B95CAE370B0582C160B8DC6E370B6CE606DE4C9988A351A0CC441;
defparam spx9_inst_0.INIT_RAM_08 = 288'h891C39B4C95CAED9AEF70BC1E10F853ADE72AAEDB2D768AA4FA32F57238DC4E371BDA111;
defparam spx9_inst_0.INIT_RAM_09 = 288'h8DB6932BA6D3EDF6BA4CA64F0582B8DFEDF5FB7DBEDF6FB75BABB4CA6D6E974BA5D2E974;
defparam spx9_inst_0.INIT_RAM_0A = 288'h4CAE5B4DA7D369B4DA6D3E9F6FB7D36972580B058B0B95CA64F0BA6D2E532583C26172FB;
defparam spx9_inst_0.INIT_RAM_0B = 288'hA9E536BB5DAFD86E37FB7D7ABD4DA757ABD5EAFD82C573C0DC2DF60B058B0993C1E132B9;
defparam spx9_inst_0.INIT_RAM_0C = 288'h41A0D06834120B2F97CB6D76D95BA5D2E93389C49E4F289CCE673389C4E26F258B45E533;
defparam spx9_inst_0.INIT_RAM_0D = 288'h0B05BEC160B0DC6E371B7D6E4AEF5519C8C451988824131189048341A8D46A351A8D46A3;
defparam spx9_inst_0.INIT_RAM_0E = 288'h28A4AABF7FBF5F6F968A94F22EF471389C6E57D4BA9F5DA54A6594FA8582DF62B9DCAE17;
defparam spx9_inst_0.INIT_RAM_0F = 288'h1BFD82C160B85FEDD6FB7DBEDB5BA5CEE973A9DCE24B0076B6D98DF70BCE291489402010;
defparam spx9_inst_0.INIT_RAM_10 = 288'h6D2E53016EA858F0782C1E172B95CAE4F0984CAE5F4FA5C9E1B4FB8DBEDB4993C1E0B058;
defparam spx9_inst_0.INIT_RAM_11 = 288'hDAED76BD5FB0582C371B8D82C371B95CF0993C26132B96D369F51B7D369F4FA7D3EDF4DA;
defparam spx9_inst_0.INIT_RAM_12 = 288'hBA552693399CCE67137934962B17944E24D158B4A6753A9D4EE994EAFD82C16FAFD7ABB4;
defparam spx9_inst_0.INIT_RAM_13 = 288'h15E224CE45198882413120906A351A8D46A351A8D46A341A0D06834165EED75CAED72B74;
defparam spx9_inst_0.INIT_RAM_14 = 288'h37138DCF0C9FD7AB7378AC1E353CA6D36BF61B95C6E16FB7DBEDF60B05C6E370B7D726EF;
defparam spx9_inst_0.INIT_RAM_15 = 288'hBA5CEA75399BC5202E0703CA0D29A6572B749A4522955CB7DC6E17FBFDFAF566A84EA0AE;
defparam spx9_inst_0.INIT_RAM_16 = 288'h7D36972B95CB69F4B94C36A36FB6DB68F2583C160AE370B85C2E370BF57EC371BFDB6B73;
defparam spx9_inst_0.INIT_RAM_17 = 288'h1B9E172994CAE5B4FA7DBEE371B7DBEDF4FA7D36974B94CA606FF6FB0DCAE572C26572DA;
defparam spx9_inst_0.INIT_RAM_18 = 288'h58B45E4F299D4EE974A9D4EA794DA757ABF5FAFD7ABD5EAF57EBF60B0582C161B0582C36;
defparam spx9_inst_0.INIT_RAM_19 = 288'h51A8D46A351A8D46A351A8D4683DBE5B2D95BA5D2A954A9CCE673399CCE6713793452290;
defparam spx9_inst_0.INIT_RAM_1A = 288'h995CF6BF60B0582C16FB75BEDF60B05C2C160B05B693146FAA8EE43110482624120D46A3;
defparam spx9_inst_0.INIT_RAM_1B = 288'h1C16070170B85C2E381C0E02E170BF5EECD509ECAA31057A39DF52B9D4A22B037A3DA0F1;
defparam spx9_inst_0.INIT_RAM_1C = 288'h5D1E06E782C0DC6E370B85C6E16EA858B017EAED32994B9DCEE73278A40DE90794D36A17;
defparam spx9_inst_0.INIT_RAM_1D = 288'h7DB69B4DA5D2E532984C9E0AE160B0DC6E373C265B51B7D36972B96D3E9B4B96D3E9B4DA;
defparam spx9_inst_0.INIT_RAM_1E = 288'hCA6D3ABF6FB7D7ABD5EAFD7EA160B7D82C160B0586E372C2E572994CAE5B4FB7DBEE36FB;
defparam spx9_inst_0.INIT_RAM_1F = 288'hCB656EB74BA5D2E995CAE572B95BA552A933893492270482C5E533A9DD32994A9D4EE794;
defparam spx9_inst_0.INIT_RAM_20 = 288'h0B0582C160B05BEB926782ECEC431104826241A8D46A351A8D46A351A8D46A351A8D47B7;
defparam spx9_inst_0.INIT_RAM_21 = 288'hFBD58E7F2E9F4F675177B3D5E8F47A3C9E4F47AC160D0995CF29B4FB0D86E16FB7DBEDF6;
defparam spx9_inst_0.INIT_RAM_22 = 288'h1B963ABB5DAED76974B9DCEA71268B46A7B50B96132B95D2E974B94CA64F2581C0DC6E17;
defparam spx9_inst_0.INIT_RAM_23 = 288'h1B8582C573C2E5F4FA6D2E532DA7D36972B95CAE572B93C0DCB0581B8DC6E171B8DC2C16;
defparam spx9_inst_0.INIT_RAM_24 = 288'h0B0582C160B0DC6E575CB6974994CAE5B4DA6D3EDF6FA5CAE572994C9E130B95C9E0B057;
defparam spx9_inst_0.INIT_RAM_25 = 288'hCADD2A95499BC9224F27A41A313BA6576BB4CA5D32794CA6D3EA16FAFD7ABD5EAFD42C16;
defparam spx9_inst_0.INIT_RAM_26 = 288'h21104C48341A8D46A351A8D46A351A8D46A351A8EEB55AAD56A975CAED7ADD6FB7DFEDB6;
defparam spx9_inst_0.INIT_RAM_27 = 288'h27138DED0894CA22F168446E7F5FB0586E370B7D82C170BFDBEC160B05BEB93778AE8EA4;
defparam spx9_inst_0.INIT_RAM_28 = 288'hB9FD4AE995CB69B4FA7D3E9B4DA5D264F2582C16071F7BB24FA3B1E97D3E99398B3D1C6E;
defparam spx9_inst_0.INIT_RAM_29 = 288'h4C160F0783C1E0F0581B8DC6E371B8DC6E370B85C6E580BF57ABF5FB7572994DA5CE6532;
defparam spx9_inst_0.INIT_RAM_2A = 288'h4CAE5B4DA6D369B4994CAE5B4993C1E132994C26132580B0586E574C2E572B95CA6572B9;
defparam spx9_inst_0.INIT_RAM_2B = 288'hA9E536BD5DA6532794CA6D3EA160B7D7ABF50B05BEC160B0582C372B95CB0996D3697299;
defparam spx9_inst_0.INIT_RAM_2C = 288'h51A8D46A351C5228F47A34E2733A9D52E995CAE572B95CAE572B7499AC49E2E179C1A333;
defparam spx9_inst_0.INIT_RAM_2D = 288'hDA058AE371B85C2E17FB7DBEDF60B05BEBB4989B710E431189048351A8D46A351A8D46A3;
defparam spx9_inst_0.INIT_RAM_2E = 288'h5D264F2793C16031B79AA5027B1C974FE9D4C94C59E6E271B9A111994462352C9E532973;
defparam spx9_inst_0.INIT_RAM_2F = 288'h1B8DC2E160B960B017FB7D82E37FB6D769B5CA5CF29D51BA6172DA6D3E9F4FA7D3E9B4DA;
defparam spx9_inst_0.INIT_RAM_30 = 288'h4C26572994CAE532580B8586E784CA6572B94CAE572782B95CAE571B8DCAE571B8DC6E37;
defparam spx9_inst_0.INIT_RAM_31 = 288'h0B7DBEC160B0582C160B0586E583C26174DA6D2E572994CAE974BA5D2E8F0784CB653278;
defparam spx9_inst_0.INIT_RAM_32 = 288'hCADD2E954AA552A974BA5D2E974A9C49A290482C5E333BA6D7ABD5DA6532994CA757EC16;
defparam spx9_inst_0.INIT_RAM_33 = 288'hFB0582DF5B9BBC598872A8D04A351A8D46A351A8D46A351A8D46A38AC566B358A5532B95;
defparam spx9_inst_0.INIT_RAM_34 = 288'hA8E4BA7F4D9D49E08E372BDE111995CFABF6EADCE2332DA0586E371B8DC2FF6FB7DBEDF6;
defparam spx9_inst_0.INIT_RAM_35 = 288'hEAF57ABB4DA7542C574C2E572D96D3E9F4FA7D3E9B4DA5D26532993C16031B7AB257A551;
defparam spx9_inst_0.INIT_RAM_36 = 288'h4CB69B4B95CAE530572B9606E160B0DCB0570B85C2E170B85FEC372C1606E161B9606FF6;
defparam spx9_inst_0.INIT_RAM_37 = 288'h4CB69B4DA5CAE4F0784CA6532994C960B0995CA60F0994CAE532784CA64F0571B95CB078;
defparam spx9_inst_0.INIT_RAM_38 = 288'hBA652E93399C4A6774CA6D3ABD5DA6D369B4DA7D7EC160B0582C160B0DC6E160B0DCB078;
defparam spx9_inst_0.INIT_RAM_39 = 288'h51A8D46A351A8D46A351A8D47159AD566B149A556A93389C4E273399CCE6733A9D52E974;
defparam spx9_inst_0.INIT_RAM_3A = 288'hEA0582DD5CA445A132DA7D42C371B85C2E170B85C2E170B8DC6E37EAD499E0BD4D19CAC4;
defparam spx9_inst_0.INIT_RAM_3B = 288'h5CB65B4DA6D3E9F4DA5D2E572993C96031977B153653077C4325D4D9DCA22AF57B3DE152;
defparam spx9_inst_0.INIT_RAM_3C = 288'h1B95CAE170B05FEDF6FB05CB0582C0DC6E582C05BABD5EAF57ABD5FA8586E573C26130B9;
defparam spx9_inst_0.INIT_RAM_3D = 288'h2C1E132B93C1E0F0983C1E0F0783C1E0F0572C1E0F0B97D36972DA6D264AE372C0DFEC16;
defparam spx9_inst_0.INIT_RAM_3E = 288'hEAED369B5EAFD42C160B0582C372B8DC2E160B960F0786D369B4BA4C9E0B0782B960F078;
defparam spx9_inst_0.INIT_RAM_3F = 288'h8A34CE45239248A07058C4E673399CCE271389CCEA774DAF5BABB5DAE532994CA757ABD5;

SPX9 spx9_inst_1 (
    .DO({spx9_inst_1_dout_w[26:0],spx9_inst_1_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_1}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_1.READ_MODE = 1'b0;
defparam spx9_inst_1.WRITE_MODE = 2'b00;
defparam spx9_inst_1.BIT_WIDTH = 9;
defparam spx9_inst_1.BLK_SEL = 3'b001;
defparam spx9_inst_1.RESET_MODE = "SYNC";
defparam spx9_inst_1.INIT_RAM_00 = 288'h1B85C6E571BFDBEC171B8DCAE170B757271136F264CE451A8D46A351A8D46A351A8DEB15;
defparam spx9_inst_1.INIT_RAM_01 = 288'h2C0636F375A953A75167B3E2152D9ED3273167ABE2393DA652E73268341E311996502C37;
defparam spx9_inst_1.INIT_RAM_02 = 288'h1B9606E17FB7DBEBF5EAF57EA160B0D86E774C1E0F0784C2E5B2DA7D3E9F4DA5D2E53279;
defparam spx9_inst_1.INIT_RAM_03 = 288'h3C1E0AE783C1E132B95CAE5F4FA4C8DC6E370B7D42DF6FB05C2C170B85BEDF60B8DCB037;
defparam spx9_inst_1.INIT_RAM_04 = 288'h2B85FEDF61B960F0DA6D369B4BA3C15C6E160B8DCB0784CA6532782C160B0572C1E0B058;
defparam spx9_inst_1.INIT_RAM_05 = 288'h89B4962D2AA5D2A93389DD3ABF6EAF5769B4DA757ABD5EAED3ABD5FB7D82C361B8DC6E57;
defparam spx9_inst_1.INIT_RAM_06 = 288'h0BFDBABB4A923B53056228D46A351A8D46A351BD5A87409643E2937A4CEA754AA5526733;
defparam spx9_inst_1.INIT_RAM_07 = 288'hC9F53A993A8CC6231188BC5E2D088DCF6994DA757EC160B85C6E17FB7DBEDF60B85C2E37;
defparam spx9_inst_1.INIT_RAM_08 = 288'h0B0D8AE782B95CAE784C2E5B2D96D3E9F4DA5CA64F038FC6DEAF165B0D3271157A395F31;
defparam spx9_inst_1.INIT_RAM_09 = 288'h1B8DC6E16FB7DBABD5EAFD82E17FB757EC370B8DCB0582C0DC2E160B05BEDF5FAFD7EC16;
defparam spx9_inst_1.INIT_RAM_0A = 288'h2B85BEDF6FB05CB0994C1E06E160B0DC6E784C0DC2DF60B0DCF0783C26572B95CBE9B498;
defparam spx9_inst_1.INIT_RAM_0B = 288'hDA6D369B4DA757ABD5DA6D3ABF60B0582C572B95CAE570BFD7EC372B9E1B4DA6D3697278;
defparam spx9_inst_1.INIT_RAM_0C = 288'h51A8D46A32A0CC27F2F8A4E6B75AA552673379345229158AC5A513BA656E954BA6536BB5;
defparam spx9_inst_1.INIT_RAM_0D = 288'hFA8D82DD5DA5CF29D5FB0582FF6FB7DBEDD6EAFD82E170B8DC6E16C9B3C176772B1146A3;
defparam spx9_inst_1.INIT_RAM_0E = 288'h6D3E9B2B94C9E071F7DBE5EEEF63AFD2E4F1479B91EF0B96CFA9D4C9CC59EAF57B41E173;
defparam spx9_inst_1.INIT_RAM_0F = 288'hDAF582E161B960F0571B8DC6E370B7DBEBF5FAFD42C161B15CEE572B95CAE785CAE572B9;
defparam spx9_inst_1.INIT_RAM_10 = 288'h0B0DCF0780BED76BF50B15CF0984C2E572DA6D2E4AE161B85BEDF6FAF5769B4EB7D82DF6;
defparam spx9_inst_1.INIT_RAM_11 = 288'h0B058AE783C0DC6E16FAFD82C573C2E9B4DA6D2E4F0580B757ABD5FB0DCF0781BFDBABF6;
defparam spx9_inst_1.INIT_RAM_12 = 288'h79AC5204F077B41C5058B4A2554CAED72B74BA5D2E774CA65329B4EAF57EBD5DAFD42C16;
defparam spx9_inst_1.INIT_RAM_13 = 288'h0B7DBABB5FB05C2E171B8DC6E37EACC4DBC99339188C451A8D47D3F98CCE6B39A5D72B54;
defparam spx9_inst_1.INIT_RAM_14 = 288'h0A64E651178AC0DE8E7864BA9F4D9CC620F0783C2E6151B05B6B5358342A5D50B05C2FF6;
defparam spx9_inst_1.INIT_RAM_15 = 288'hFB7D7ABD5FA8582C361B95C6E371B95CF0984CA6572D96CAE572B93C0E3EFD7EBEDE6EB6;
defparam spx9_inst_1.INIT_RAM_16 = 288'h6CBE9B4D93C0DBEDF6EAF57ABD5DA6D369D5FB7DBEDB5DAF57EC372C160AE582C1606E16;
defparam spx9_inst_1.INIT_RAM_17 = 288'h5CB69F4DA4C9E0B017EAED76BD50B0DC6E16DAED3AA161B95CAFF6DAED7EC161B15CF098;
defparam spx9_inst_1.INIT_RAM_18 = 288'hA9D52E994BA4CEA794CA65369D5FB05BEDF5FB0582C371B8DCB0581B85C2DF60B0586E78;
defparam spx9_inst_1.INIT_RAM_19 = 288'hFAED2202CB3C1588A351A8FE6747ACD66B55AAD5628B2287BB9BADE6FB85C7058BCA6733;
defparam spx9_inst_1.INIT_RAM_1A = 288'hFA7D3673167BC2E793A93C5608F47BC6A7F50B8DC6E370BFDBEDF6FB05C2C160B05C6E16;
defparam spx9_inst_1.INIT_RAM_1B = 288'h2B960F0784CA6572B95CAE532781C05FEFF7EC5DDAC14D9DCEA75399445E2D078442A5B3;
defparam spx9_inst_1.INIT_RAM_1C = 288'hDA757ABD6FB75B6B94CAFD86E371B960F0993C05C2DF6EAF57ABD5FA8582C361B0D82C36;
defparam spx9_inst_1.INIT_RAM_1D = 288'h0B05BEBB4CA757EC372B95FADF60B0D82C161B9E130FA7D2E530570B757AB94B9DCF2794;
defparam spx9_inst_1.INIT_RAM_1E = 288'h0B7DBEC161B8DCAE782C160AE370B0DC6FD5FB15CF0995CB69F4994C9E02DD5EAF576BF6;
defparam spx9_inst_1.INIT_RAM_1F = 288'hAAC51A8B43A14CA451281C120B158AC5207038241A31299D4EA753A9D4EE794B9E53AA16;
defparam spx9_inst_1.INIT_RAM_20 = 288'h8954AE793DA7DBEDF60B0DC2E160B7DBADD6EB7DBEC170B756628E05D1DC8A351B56AD96;
defparam spx9_inst_1.INIT_RAM_21 = 288'h0B85C31F8BBBD8ABF4C9DCEE753A9D4E651178BC263B30A8D7A97298CC9E0AF47A4160F1;
defparam spx9_inst_1.INIT_RAM_22 = 288'h2C1E0B0580B85FEDD5EAF57ABD5FB0586C360B0586C372B95CB0984CA6572B95CA64F038;
defparam spx9_inst_1.INIT_RAM_23 = 288'h1B8D86C373C1E1F4FA5CA60AE16EAF572752A95CF2794DAED7ABD5DAE52E974EAFD82C37;
defparam spx9_inst_1.INIT_RAM_24 = 288'h0B05BABF60B96132B96D3E932993C0DFABB5DAED7EBF5EAF5329B4DA7546E782BE53EC37;
defparam spx9_inst_1.INIT_RAM_25 = 288'h79349A2B13824162F28944A6753B9E532994CA7542C370B0586E572B960F0993C15CAE17;
defparam spx9_inst_1.INIT_RAM_26 = 288'hEB6D76BD6EB7D82E170B756E71036EA64AC4CB65AAAD419048263319948E27148AC5A2F2;
defparam spx9_inst_1.INIT_RAM_27 = 288'hB9DCEE75378B41E192FA0542BD4B9B3CDC8F683C6A573A9CC9E331B9DD36A161B8DC2DD6;
defparam spx9_inst_1.INIT_RAM_28 = 288'h0B0582C160B0D86C371B95CF0984CA6532B94C9E0B0381C0E3F1978B2546BD4B9D4EA773;
defparam spx9_inst_1.INIT_RAM_29 = 288'hDA5CEA553B9E4F29B4DAED76BB5CA5D2A7B4DAFD86E583C1606E370B7DBABB5DA6D7ABF6;
defparam spx9_inst_1.INIT_RAM_2A = 288'h1BF5769B4DA6D76994CA65329B4EA95CF037DA858AE571B95CAE784C3E9F4B94C15C2DD5;
defparam spx9_inst_1.INIT_RAM_2B = 288'hCA6D369B4EA8586E371B8DCF0782C1E172B93C9E06E16FB7DBEDF61BA6132B96D264F078;
defparam spx9_inst_1.INIT_RAM_2C = 288'h577AACFB6AAAD02550B87C8A673391C8E270381C1209168BC9E4D158AC5E4F27944A6573;
defparam spx9_inst_1.INIT_RAM_2D = 288'hA8B3D9EF088D4AE7539944A22F0785CFEC371BFDBABD6EB7DBEDD6FB7DFEDF6EB7576952;
defparam spx9_inst_1.INIT_RAM_2E = 288'h4CA6572993C960B0581C05F6F577B1D7E993B9DCEA753B9E532953893415F10C98D46DF4;
defparam spx9_inst_1.INIT_RAM_2F = 288'hBA54F2994EA85CB0994C95C2FD5DA6532994DAF57EC160B7DBEA160B7D82C371B960F078;
defparam spx9_inst_1.INIT_RAM_30 = 288'h2B95C2C162B9DC6E163C260F0997D3E8F0782B85B6B94A9D4EE773CA6D32994CA6536B95;
defparam spx9_inst_1.INIT_RAM_31 = 288'h3C1E574DA3C15C2DF60BFDBEC373C1E132B93C15C6E37EAE5329B4CA5CEE793CA65329D5;
defparam spx9_inst_1.INIT_RAM_32 = 288'h49244E04F077BBDC0E282C5A4F27944A25128944AA794DA75769B4EA8582C161B9E13078;
defparam spx9_inst_1.INIT_RAM_33 = 288'h997546E572B8DC2DD6DAF5BADF6FB7D82FF6EB7576973882362AB409DC61F901924D2692;
defparam spx9_inst_1.INIT_RAM_34 = 288'h5B0D7A993B9D4EA753A9D4EA75399445E2D098F506A35EA5C9E0AF573C222F1582C1A0B0;
defparam spx9_inst_1.INIT_RAM_35 = 288'hCA5CF29D5FAFDBEDF6FA8582C160B0582C161B95CF0994CA6532782C160B0580BF5EEF36;
defparam spx9_inst_1.INIT_RAM_36 = 288'h5C95CAE983C7DAE753A9DCEA773DA6D72974CA7572B74A9D4EE9D51B96132780BED72994;
defparam spx9_inst_1.INIT_RAM_37 = 288'h2C1E132581B8DC6FB5B9DCEE753A954EE794DA6D368370B754AE572B8DC2C574C26532DA;
defparam spx9_inst_1.INIT_RAM_38 = 288'h58BCA25329954F29D5DA65369D5FAFD82C162C26574B95CAE572992C0DC2E161B8DCAE57;
defparam spx9_inst_1.INIT_RAM_39 = 288'hDAFDBADD6EB75BABB4B914C27B2B8E43E252291C8E471389405FEED66339BEE078BC5E50;
defparam spx9_inst_1.INIT_RAM_3A = 288'hA9CC9E2D098E4C2A15FADC99E8E4733D5E6E3734265D40B05BEBF61B85FADB5DAED7ABD5;
defparam spx9_inst_1.INIT_RAM_3B = 288'h0B7DBEC171B96132994CA64F0783C1607017EBE5EAEF64A8532752A94CA25129954EE773;
defparam spx9_inst_1.INIT_RAM_3C = 288'hDA652E9B4EB652A733995CFAA172B9606FF6CA652E973BA6D7EBF60B0582C160B05C6E37;
defparam spx9_inst_1.INIT_RAM_3D = 288'hB9E5369B4CA6D02DF5EA9E0AE371B8DCF0B95CA6172982B8DCF0991BE52A753994CAE794;
defparam spx9_inst_1.INIT_RAM_3E = 288'hEAFD7EC373C2E9B4DA6D36972782C0DC6E371B960AE583C1E0B0160B0DFAB73A95CEA552;
defparam spx9_inst_1.INIT_RAM_3F = 288'hD8F442452190C422312813C1DCDC6633198CB652ED9EE483462532A9E53ABB5DA65369B5;

SPX9 spx9_inst_2 (
    .DO({spx9_inst_2_dout_w[26:0],spx9_inst_2_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_2}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_2.READ_MODE = 1'b0;
defparam spx9_inst_2.WRITE_MODE = 2'b00;
defparam spx9_inst_2.BIT_WIDTH = 9;
defparam spx9_inst_2.BLK_SEL = 3'b001;
defparam spx9_inst_2.RESET_MODE = "SYNC";
defparam spx9_inst_2.INIT_RAM_00 = 288'h57A389A6E88ED0AE770B54AA5B4FB7DBADB5CAE532994DAED7ADF60B7DBEBD5E96CB63B1;
defparam spx9_inst_2.INIT_RAM_01 = 288'h2C0DC2FF7EBE5E6EB61AECEE5328944A6573CA652E753A9CCA24F1785CB69D4DA64EA2F0;
defparam spx9_inst_2.INIT_RAM_02 = 288'h1B85FEDD5CA5D2E994EAFDBEC161B8DC6E371B8DC6E16FB7D82C372C1E132994CA653299;
defparam spx9_inst_2.INIT_RAM_03 = 288'h2BA6172B93C1E0AE371B9E13057DA5CEA712894CAE794B9DD36BD5CA4CE2512A9ED7EC37;
defparam spx9_inst_2.INIT_RAM_04 = 288'h1B8DC6E372B960B0582C0DFEDD50B756E752A94CAA794DA75369B4EA7D7ABF53B95C6E57;
defparam spx9_inst_2.INIT_RAM_05 = 288'hC652E972A8542A97EE483C66573CA757ABB5DA65369B5EAFD42C373CAE9B4FA6D2E53258;
defparam spx9_inst_2.INIT_RAM_06 = 288'hEAFDBAD94BA65329B5DAF57EDF6EB757ED91D8F4BA390D87C465F1E8EC7E251489C05FCD;
defparam spx9_inst_2.INIT_RAM_07 = 288'hB9E532994B9D4EA73299D4EE75388BC1E1720A857271057239A1730B0D86DD599341E373;
defparam spx9_inst_2.INIT_RAM_08 = 288'h2B8DC6E370BFDBEDF6FB7D82E382C1E0F2794CAE532581B8DC2E17DBD5DAC54D9DCA6532;
defparam spx9_inst_2.INIT_RAM_09 = 288'hB9D4E2512894CB2973BA6532994A9C4A2553CA758AE572B8DC2DD5DAED7ABF6FB7D86E57;
defparam spx9_inst_2.INIT_RAM_0A = 288'hEAED2A5119954F2794FAF5769D5EAF542C572B95CAE574C2E572572B8DC6C373C1E06D94;
defparam spx9_inst_2.INIT_RAM_0B = 288'hEAFD7EBD5DA65369B5EAFD82E584CB69B4DA5C9606E171B85C2E372C160AE371BFD76BD5;
defparam spx9_inst_2.INIT_RAM_0C = 288'hEA85B23D2E96469FD1097CB6371C8F44E2D2692401DACC663319ADD6E339A6F78D4F29B4;
defparam spx9_inst_2.INIT_RAM_0D = 288'h89341E172D9F53E9D4D9E4EE772A94C622D0582C1E312A9E53AA160B7DBABD6EAE536BB5;
defparam spx9_inst_2.INIT_RAM_0E = 288'h2C160F2BA5D264F0582C16071D7BBB54275188446A573CA5D2E7328944A6553CA6D32973;
defparam spx9_inst_2.INIT_RAM_0F = 288'h793462574FB1E0F0571B8DC2C171B85C6E372B8DC6E572B85BEDD5DAED76BD5FB0586E38;
defparam spx9_inst_2.INIT_RAM_10 = 288'hEAFD8EE783C15CEE985C9E02C161B95C6E371BFDB6994A9C4A24F1895D2A753BA5D2E953;
defparam spx9_inst_2.INIT_RAM_11 = 288'h5CB69F4B92C05BEDD5EB7D82C371B8DC6E17FAED329B5DA54DE311B9E5327F60B75769D5;
defparam spx9_inst_2.INIT_RAM_12 = 288'hA8740E2B1481BC9E4F379C1209048241A312CA6D3ABD5EAFD7EBD5DA6D36BD5FA8586E78;
defparam spx9_inst_2.INIT_RAM_13 = 288'h4723D5EB0482C1A132B9ED7EC160B0582DD5BA5D32BD5EAEC7E5D2C8F4423F2D9646E350;
defparam spx9_inst_2.INIT_RAM_14 = 288'h3A645DEEF784C6A552994CA65129954EE794DA6D36B94A9CCAA552B9750AC761B6D262AF;
defparam spx9_inst_2.INIT_RAM_15 = 288'h1B8DCAE571B85BEDF6EAED72973A9DD329D5FB05C2E372C1E532994C9E4F0783C0E3AF56;
defparam spx9_inst_2.INIT_RAM_16 = 288'h1B8DC2DF5EAF57295399449E312B9D4EA753BA55266F158346A7F62C15CAE582C15CB078;
defparam spx9_inst_2.INIT_RAM_17 = 288'h1B8DC2DD5CA5CF2994B9C462373CA5CC2C37FADCF6BF50B1DCEE572B9DD30B94C0D82C36;
defparam spx9_inst_2.INIT_RAM_18 = 288'hA9D4EA794EAFD7EBF5FA85BEBD5DA6D36BD5FB058B0795CAE93257FB6D32994EAFD82C17;
defparam spx9_inst_2.INIT_RAM_19 = 288'h2B95C2DD5CA6536BB5C8EC763B1F8F4763B2C8DC6A150C80C0E07038241A2F17944AA753;
defparam spx9_inst_2.INIT_RAM_1A = 288'hB9DCF2994CA7576BB5DA652A711A9054AC560AE4E62CF47ABD60B068446E794DA5CEE7D5;
defparam spx9_inst_2.INIT_RAM_1B = 288'h995D36BD5FB05C2E382C1E4F2783C1E0F0781C7DE6A32A843DDEEF783C1E0F088CCA6553;
defparam spx9_inst_2.INIT_RAM_1C = 288'h99CCE675399BC960906854FEC160B8DCF0783C1E0AE571B85C2FF6DADD2E753A9C4A2512;
defparam spx9_inst_2.INIT_RAM_1D = 288'hB98586DD5B9F57EC363C15C2C373C2E1B2B93B8582C160B7D7ABD5FB6D6A73278B45E353;
defparam spx9_inst_2.INIT_RAM_1E = 288'hDA6D36BD5FB0DCB0794C9E02DB5B9D4EE794EAFDBEC161B85F6973B9D4F29949944AE794;
defparam spx9_inst_2.INIT_RAM_1F = 288'hA85C765B2D8EC7A3F1289C49E4F382C5A312A9DCF2994CA65369F50B0582DF6FB7D7ABB4;
defparam spx9_inst_2.INIT_RAM_20 = 288'h98D4B27F41B7D6E4F057ABDA111A9653ABD5A934222164C2606FD5DAED76B70B8643A190;
defparam spx9_inst_2.INIT_RAM_21 = 288'h3C1E0B038EBC54A591A83BD9EAF57A391CD09954EE773A9DCEE773CA65329D5EAF572912;
defparam spx9_inst_2.INIT_RAM_22 = 288'h1B9E172B94C8DC6E16FB756E91258B4560B0582C1E333CA6D7ABD6FB05C6E381C160B058;
defparam spx9_inst_2.INIT_RAM_23 = 288'h4C2E5B2B91BFD42DF5EAED3AA16DAD4E24D15834625128944A24F2581BCDED1A9F57ABF6;
defparam spx9_inst_2.INIT_RAM_24 = 288'h994CA6774DAF57EDF60B6526532995D329329954F2994FB05BAB94FA858AEB92B8DCAE98;
defparam spx9_inst_2.INIT_RAM_25 = 288'h0713CE0D1894CAE794DA753ABF50B0582DF5EAF57ABD5DA6D3ABF60B16132791BF572953;
defparam spx9_inst_2.INIT_RAM_26 = 288'hB9ED3EDB5C9E53EA162B9DC6FF5DAED6A170C853DDD0FB86CBE432299CD26B3591C05DED;
defparam spx9_inst_2.INIT_RAM_27 = 288'h271B95EF078446A552B9E4EE753B9ED3ABF5DAE52E73388BC223B40AFD7693167A399F52;
defparam spx9_inst_2.INIT_RAM_28 = 288'h171BD61129954EE794EAFDBEDF60B05C2E371B8DC6E381C0E02FB68A94B210F67ABD1E6E;
defparam spx9_inst_2.INIT_RAM_29 = 288'h99BC5609058345A2D168B45202F07139A353DA6D7EC373CAE532580BFDB2B53892C49E2E;
defparam spx9_inst_2.INIT_RAM_2A = 288'hB9DCEA732A9E5369D50B05BEA161B95CF0572BA6170B96CB657216FA85BEDB4CA757EDB5;
defparam spx9_inst_2.INIT_RAM_2B = 288'h0B0D82DD5EAFD7EDF5EAFD82E371B9E13258FB652651278BC66594DAF57ABD5CA4CA6532;
defparam spx9_inst_2.INIT_RAM_2C = 288'h1BD42A14F772B59D0FC8FC8E6D47A45228F35893C1C0E27A41A312A9E4F69D4EAFD7EBF5;
defparam spx9_inst_2.INIT_RAM_2D = 288'hCA6536B94BA652E97499C4AA572EA0546BB38833DE111A9F546C572B8DBEDD5EA8582C36;
defparam spx9_inst_2.INIT_RAM_2E = 288'h0B05C2E171B8DC70381BFDF6D3529DC1DEAF47238DC4E372BD5E8E57C466573B9D4A6553;
defparam spx9_inst_2.INIT_RAM_2F = 288'h07346A7B5EB7D82E783C0DFEDB5BA4CDE290278B85C6F68D4F69D5DAED7ABD5FB0582C16;
defparam spx9_inst_2.INIT_RAM_30 = 288'h1B8D8AE773C261B2D94C1DFABD50B7D6E953DAF5B2912481BC9E6F481BD20903803B9BAC;
defparam spx9_inst_2.INIT_RAM_31 = 288'h3C1E0F037DA4C9E2D068BC6A794DAED769739944A2552B9D4EA552B9ED7AA161BFDBEC16;
defparam spx9_inst_2.INIT_RAM_32 = 288'hAAD52A913689BC9E907954EE794DA753ABF5FAFD7EBF50B05BEBF5FA8582C161B95CF058;
defparam spx9_inst_2.INIT_RAM_33 = 288'hEA25CEDF4B94419EF0B9058EE983C0DAE6F0B9FD4AE98A853E1ECE673BA5F91F924DE934;
defparam spx9_inst_2.INIT_RAM_34 = 288'hB833D5C8E47238DC8E57A38DC8E67C466552994CA6552A9DD2E974CA6536BD6EB5D22311;
defparam spx9_inst_2.INIT_RAM_35 = 288'h68AC0DE2E171BDE373EA8D86C160B7D82C160B05BEDF6FB7DC2E371C160B0380BF5EAC73;
defparam spx9_inst_2.INIT_RAM_36 = 288'hEADCEA794DADD1A24F270B85C4F170B85E0ED65AED7EE78DD36BF6EB0586FF6DADD224F2;
defparam spx9_inst_2.INIT_RAM_37 = 288'hCA5CEA7539944A6553A9CCA6573DAED7EC16EAF57EA160B1E130774C36572781B6D369F5;
defparam spx9_inst_2.INIT_RAM_38 = 288'hEAFD7EBF5FAFDBEBF5EAFD7EC160B0DCB0782C1E0F2782C1606FD5A93411E905844AE7B4;
defparam spx9_inst_2.INIT_RAM_39 = 288'hFADCDE2D0896D02D90C8642DF90E8848A4936A452AB75CAED72B54893CA6794EAFD7EBD5;
defparam spx9_inst_2.INIT_RAM_3A = 288'h783C22352A94CA6573BA54EA794BA657EC170BED624F0D98546C560ADC95CAE98E53EA16;
defparam spx9_inst_2.INIT_RAM_3B = 288'h1B0582C160B7DBEDF60B85C2E382C160B0581C5DCE750572B99EEF57A391C8E47A3D1EAF;
defparam spx9_inst_2.INIT_RAM_3C = 288'hD66B3596BA5DAC1CD1A9E536BD5EAE5266F24813C5E2EF6EB2976BF73C76A362B95CAE57;
defparam spx9_inst_2.INIT_RAM_3D = 288'hCA7542DD5EAFD82C163C260F0B96CAE4EE37FAED369B4CA5D2E974A9AC41DEDF68381DCD;
defparam spx9_inst_2.INIT_RAM_3E = 288'h1BA6532781B8DCB0581B85BAB53681BC9C6F78DD32953A9CCA65328944A2532994CAA7D5;
defparam spx9_inst_2.INIT_RAM_3F = 288'h9ADD72DB6DB6DBADF6FB75BADB5EAFD86E371B05BEBD5FAFD42C361B0DBEDD5DAFD46E37;

SPX9 spx9_inst_3 (
    .DO({spx9_inst_3_dout_w[26:0],spx9_inst_3_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_3}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_3.READ_MODE = 1'b0;
defparam spx9_inst_3.WRITE_MODE = 2'b00;
defparam spx9_inst_3.BIT_WIDTH = 9;
defparam spx9_inst_3.BLK_SEL = 3'b001;
defparam spx9_inst_3.RESET_MODE = "SYNC";
defparam spx9_inst_3.INIT_RAM_00 = 288'hBA6D7EC17FB5D2251198DCBA8561B6CE20CF784C6E75278AC11E8F58444625239249A714;
defparam spx9_inst_3.INIT_RAM_01 = 288'h2C1E4B2189B04A5EEF884C1E0AF47A3D1C4E269B95ECF57B422331783C265539944A6553;
defparam spx9_inst_3.INIT_RAM_02 = 288'h588BFDD8C95C29D288239A2562F99FD8AE784C260EE370B7D7ABD5FB7DBEDF6FB85C6E38;
defparam spx9_inst_3.INIT_RAM_03 = 288'h3B95C6DF5FAFDBAB94BA5D26712487B79BACD66B2D74BA5D2E574BD61BE6574BA5CEE933;
defparam spx9_inst_3.INIT_RAM_04 = 288'h479391ED1A9D4E651278BC6231288BC62532894CB6974DAFDBABB4DA7D42C161B15D3078;
defparam spx9_inst_3.INIT_RAM_05 = 288'h2B95CAE360B7D7EA160B0D86C372B95C2DF60B0DCAE785CAE972792C15CAE370B7572911;
defparam spx9_inst_3.INIT_RAM_06 = 288'h0AFD367305733D1E4E279BC9C4E47B4E2954BAE57ADF7FB85C2E170B85C2E170B85C2E37;
defparam spx9_inst_3.INIT_RAM_07 = 288'h57A3C9A4D372391C8E57BC1E0AF57BC665328944A6553CA75BADD6DAED6E912683C3A615;
defparam spx9_inst_3.INIT_RAM_08 = 288'h0B1E170B94C15C6DD5DA6536BD6EB75BEDF6FB85C6E582C0E3AEF509E46A1508833D1CAF;
defparam spx9_inst_3.INIT_RAM_09 = 288'hF6EB2D74AA54AE572B95CAED7ED58D4EA71278B44E1ADA5BA91227F36120723246312153;
defparam spx9_inst_3.INIT_RAM_0A = 288'h68C4A651299652E994EAF572773DA05BABF52B9E06C362B85BEA161B6D6E753A9BC9604F;
defparam spx9_inst_3.INIT_RAM_0B = 288'h2B9E0AE371B96132BA6D36972993C1606E37FB756A6B047AC1A111893C5A2B058341E2D1;
defparam spx9_inst_3.INIT_RAM_0C = 288'hBA657ADF6FB05C6E371B8E070381C0E070582C1E0F0782B8D82C161B0582C161B0D86E57;
defparam spx9_inst_3.INIT_RAM_0D = 288'h684466532A9CCEA774DADD329D50BFDB2B325834223931A9DC2B10369349C6F47A3D60F0;
defparam spx9_inst_3.INIT_RAM_0E = 288'hEAF582E170B8DC70380C75E2C7409E4620CF57A3D5ECF479B8DC8E371B8DCAF67A38DC8E;
defparam spx9_inst_3.INIT_RAM_0F = 288'h792C49E0EE6DB1D4892479B0B036138B4B0B17BCB28575CB6572781BFD72773CA6D7ABB5;
defparam spx9_inst_3.INIT_RAM_10 = 288'hEAED3EA573C0D82C16FA8582C16CA54E65125813C1DACC652A150A9552E974BB66301CD1;
defparam spx9_inst_3.INIT_RAM_11 = 288'h3C8DC6E16FB6D224B0683C5E2D05823D1E6F37A3D1E9068C4A6573CA5D329B4EADCAA593;
defparam spx9_inst_3.INIT_RAM_12 = 288'h1C160F0994CA60F0370B0586C360B0582C160B0582C372C260AE583C26572DA6D2E53299;
defparam spx9_inst_3.INIT_RAM_13 = 288'hEB6DB2B74A9BC51EF01A9DC2B114723DA0F0682C1A1B5DB7DBEDF60B8DC6E382C160B038;
defparam spx9_inst_3.INIT_RAM_14 = 288'hA8C41E0CF57B3D5E8E272395EAF371349A4D269B8DC8E57C46A794B9D4EA77399D4EE9B5;
defparam spx9_inst_3.INIT_RAM_15 = 288'hA22201F12EA961B4FA6D260AFD5A9CCAE794CA6D7ABD5FB05C2E170B8DCB0590C5DD29D2;
defparam spx9_inst_3.INIT_RAM_16 = 288'h99449E29017736D72A8542A152BB6633198CD6839204FE6DB2570A651234D2481C11C6A2;
defparam spx9_inst_3.INIT_RAM_17 = 288'h271385C0D170B89C9078CCAA753B9E5369D5B94CAA7B4DA7546C782B8582C360B7D7AB73;
defparam spx9_inst_3.INIT_RAM_18 = 288'hEAF57EBF5EAFDBEDF61B95CAE583C16132DA5CA64F2792C05C2DF6FADCDE2D078C49A28F;
defparam spx9_inst_3.INIT_RAM_19 = 288'h993411C6E57C476BD6FB7DBEC171B960B0582C0E06E372C1E132983C0DC2DF6FB7D7EBD5;
defparam spx9_inst_3.INIT_RAM_1A = 288'h479B85A2D269B89C6E47B422332B9DCE6512A9E536BB5DAED7ADF6DACCDA131EA0576993;
defparam spx9_inst_3.INIT_RAM_1B = 288'h88D4EE794CA6D76BD60B8DC6E372C1E4F239BB9D3233188C422110682BCDC6E372BD5EAF;
defparam spx9_inst_3.INIT_RAM_1C = 288'hC6EB6D9AD0703B190A549200FC6A2308826261A894227C62C76A575CB69B4981B6D264F1;
defparam spx9_inst_3.INIT_RAM_1D = 288'hA9DCF29529954B2794EA058AE570B0582DF5DAED2A732893449FEEC64AA150A95DB31BAD;
defparam spx9_inst_3.INIT_RAM_1E = 288'h1B96132994C9E0F0582B85BABD5CA4C9E2F199449604E06FB399CC068B89CD0894CAA753;
defparam spx9_inst_3.INIT_RAM_1F = 288'h3C9E4F0581C0DC6E784C260F0370B05BEDF5EAE532794DA757ABB4DA652E953BA6D7EC17;
defparam spx9_inst_3.INIT_RAM_20 = 288'hB9CCA6553CA6D72B94CAF542FF7DAD4E2531B95CFA9D4D9CC59ECF886D7AC170B8DCB078;
defparam spx9_inst_3.INIT_RAM_21 = 288'h3C9E433772A5C6631088CC662F057A3CDC6E472BD5EAF471349A4E271345A2D26A39E373;
defparam spx9_inst_3.INIT_RAM_22 = 288'h51A08C26150E161670AA058F0994C9E02D9488B41E311A95CEE974CA6D7EC171B8DC6E58;
defparam spx9_inst_3.INIT_RAM_23 = 288'hFAFD7ABB5DAD4E6712480BF9B6B854AA978CE683BDDADB64AED9ADA5B2491E6C2C918461;
defparam spx9_inst_3.INIT_RAM_24 = 288'hB9CCA2332993C4DE2DF673357CC068B8DEB0894CA6512995CEA532995CF27B4FA8DC6E16;
defparam spx9_inst_3.INIT_RAM_25 = 288'hFB7D7AB94B9D4AA573CA64EE753993C560D1895D36A161B8DCB0582B8DCB0370B6D72994;
defparam spx9_inst_3.INIT_RAM_26 = 288'hEB6D6A6B047D4BEA561AF4EE330EB7D86E582C1E0F2793C1E0B0382C1E132983C15C2C16;
defparam spx9_inst_3.INIT_RAM_27 = 288'h57A3D1E8E47ABD5E8E372391C6E168B41A2D26ABE2352A9CCA6553B9DCEE994CA6D76BB5;
defparam spx9_inst_3.INIT_RAM_28 = 288'hFAE4E64F178BC62332A9DD2E994EAFD86E371B8DC6E581C062AE54C8D46211088CC622F0;
defparam spx9_inst_3.INIT_RAM_29 = 288'hC66B7DC0F38143DD2B85429D468F3595C6C271B0D450561985032454FB9E7D52C2653057;
defparam spx9_inst_3.INIT_RAM_2A = 288'h068349CB078B41A312A954A2311B9E4F27B40B05BEBD5EAED36BD5CA4C9A270076B6D74B;
defparam spx9_inst_3.INIT_RAM_2B = 288'h5824162B1795536BD6EAF57ADD6FB0DC2DF6EADD2A773A9CCA6753893451E2EF6EAF57CC;
defparam spx9_inst_3.INIT_RAM_2C = 288'h0B8DCB0783C1E0B0371B8DCB0784CAE4F0571B7DBEBD5EAED2E753A954AA753A9D4A64F1;
defparam spx9_inst_3.INIT_RAM_2D = 288'h068B49A4E372BDA0F088C46233288CCAE794CA6D76BD6FBFDB6B5378C4725D33B2586BF6;
defparam spx9_inst_3.INIT_RAM_2E = 288'hFB05C6E371C160B0580C5DD29B2983C1E11098CC620AF47A3D5ECF683415E8E57ABD1C4D;
defparam spx9_inst_3.INIT_RAM_2F = 288'h51185450381A09046120C0C91AE58D502C785CAE46FB499445E2D078C4A6553BA5D329B5;
defparam spx9_inst_3.INIT_RAM_30 = 288'hB9DCF29F5EAED32994CA652E773892C0DFEED6E32D9ED179C122D2588BDD4A9449234B03;
defparam spx9_inst_3.INIT_RAM_31 = 288'hEAF576B95CA54E65329954E6532993C9606F06F3399EDE6034DEB047B4265529944A6552;
defparam spx9_inst_3.INIT_RAM_32 = 288'h5CA60B0370B7DBEBD5DA6532994DA6D369B4CA549E2B0482C5A4F2793C9E51299E52E974;
defparam spx9_inst_3.INIT_RAM_33 = 288'h88DCEE794CA65329B5EB75B6B53893C1E1B22AADFEDF60B8DCB0582C0DC6E171B960F099;
defparam spx9_inst_3.INIT_RAM_34 = 288'h883C1E0F0783C1A0D068341A0F06833D1EAF479B85A2D269B89C4D371B91CAF683C222F0;
defparam spx9_inst_3.INIT_RAM_35 = 288'hFB1E130982BF56A4F178B45E311994CAA773BA657ABF60B8DC6E381C0E031B77A9536530;
defparam spx9_inst_3.INIT_RAM_36 = 288'h4813F9BACC66B45EB17944E6913383A91247D2B8CC22020A8A06E3410800103246352354;
defparam spx9_inst_3.INIT_RAM_37 = 288'hA9CCDE290177B7DBCCF68B89C4E47BC6651188CCA6532A964FABD5DA6D2E793B9D4EA712;
defparam spx9_inst_3.INIT_RAM_38 = 288'hFA8582DF5DA54E24D168BC9E4B13813C9E7058B45A312994CE6733893C5E312994CA6553;
defparam spx9_inst_3.INIT_RAM_39 = 288'hA9BC19F721AFD82E371B95CAE571B8DC2E373C26532983C160AE160B7DBABD5DA6D369D5;
defparam spx9_inst_3.INIT_RAM_3A = 288'h57ABD1E6E268345A6E371349A4D168B45A6E67B41E131A954B6994A9DCF6BB5DAFDBEDB5;
defparam spx9_inst_3.INIT_RAM_3B = 288'h9954EA794DAF5BEC171B8DC2E170BF5EACB409E4A6310783C1E0D078441E0F057ABDA0D0;
defparam spx9_inst_3.INIT_RAM_3C = 288'h759238CE330904824140B09848151719556D38CCFAC574C2606FB4993C5A0D068BC66532;
defparam spx9_inst_3.INIT_RAM_3D = 288'h47BC1E2F188CCA6532A9ED369B4DA5CEE753994C9E29017F37598CE693DA554BA5D2A891;
defparam spx9_inst_3.INIT_RAM_3E = 288'hC66335BCDF70381C2E27A4120904824160F1894CAE774BA54DE4901703799CCE67B01A2E;
defparam spx9_inst_3.INIT_RAM_3F = 288'h1B8DCB0994C9E0F0582C15C6E16FB757ABD5EAF57ABF50B0D82C16FAED2A7125893FDDAD;

SPX9 spx9_inst_4 (
    .DO({spx9_inst_4_dout_w[26:0],spx9_inst_4_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_4}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_4.READ_MODE = 1'b0;
defparam spx9_inst_4.WRITE_MODE = 2'b00;
defparam spx9_inst_4.BIT_WIDTH = 9;
defparam spx9_inst_4.BLK_SEL = 3'b001;
defparam spx9_inst_4.RESET_MODE = "SYNC";
defparam spx9_inst_4.INIT_RAM_00 = 288'h06FB05A6E47BC26352996532973DA75B6B94FB0DC6FF6EACC9E1110B8DC6E371B95CAE37;
defparam spx9_inst_4.INIT_RAM_01 = 288'hDBD5969F2B8CC6211088446233198B415E8F57BC1E0CF57A3CDC2D060309A6E269389A2D;
defparam spx9_inst_4.INIT_RAM_02 = 288'h9603CE313EA8DCAE571BF56A6D058345A2D188CCA2532A9DCF29B5EB7D82E170B85FEFF7;
defparam spx9_inst_4.INIT_RAM_03 = 288'hB9D4A24F178BC5202EE6E3319CD17B4AA995BA4CCE2EAE348CC26130984826140A0A07C6;
defparam spx9_inst_4.INIT_RAM_04 = 288'h178389E9068CCEE974B9D4DE290277B3578BB5733DA2E47AC160D0A954A2532B9DCEE794;
defparam spx9_inst_4.INIT_RAM_05 = 288'hEAF57ABD5EAF5369B4EA8586E572BF56A690C62A4CE674432A152B95C2A574BB66B3DA0E;
defparam spx9_inst_4.INIT_RAM_06 = 288'hDAE52E9B5FB75BADF6EB652E6171B8DC6E371B95CAE572C1E132993C15CAE571B8DC2FF6;
defparam spx9_inst_4.INIT_RAM_07 = 288'h783C1A0D088C45E0D0682385A0C169389C2D169391C8E16FB05A6E67BC1E0F0A95CEE7D5;
defparam spx9_inst_4.INIT_RAM_08 = 288'h78C462312894CAA774CA65329B5FB7DBEC170B85C31D7BB2D3E55088442635188B41E110;
defparam spx9_inst_4.INIT_RAM_09 = 288'h99E576B758994195855128544A240984C2618189EDA30594CFAA574C1E06FB4993C5E2F1;
defparam spx9_inst_4.INIT_RAM_0A = 288'h17733174AC5F305A4E47A3DA13299445E3118954EE732893C5E2F168A409FEEC65B3DC90;
defparam spx9_inst_4.INIT_RAM_0B = 288'h3C0DEE870959A38B64C2E97CC060309C8E68443A6556BB663319CD3844AE774B9CCDE290;
defparam spx9_inst_4.INIT_RAM_0C = 288'h1B8DC6E573C1E0F0984CA64F0370B0D86E371B8DC2DD5DA6D3ABF5FAF572773DA858AE78;
defparam spx9_inst_4.INIT_RAM_0D = 288'h472BD5E6E372391C4D060309AAF67ABD9EF088D4B2994DA6D7ABD6EAED7EDF6EB6D7ADF6;
defparam spx9_inst_4.INIT_RAM_0E = 288'hFB05C2E371C0E031764A6C620CF67BC220F068341A0F088BC1A0F0783415ED0478B45A4D;
defparam spx9_inst_4.INIT_RAM_0F = 288'h60D904EEAC6941A554EA95CF037EAE52651188C4A2311894462532A9DCEE974BA6536BD6;
defparam spx9_inst_4.INIT_RAM_10 = 288'h78BC5A0F19954EA71168B45E2B0481BC1D8CC60396354DAF5AEB1317A2688A1612890261;
defparam spx9_inst_4.INIT_RAM_11 = 288'h91C8E8964D28188E68442A1934B27C4AE974A9CCDE29006E2ED56AE60345C6E47BC66511;
defparam spx9_inst_4.INIT_RAM_12 = 288'h0B0586E160B05BABB4DA757ABF5FAF572994DAFD8AE983C0DEE870B6328514450A058503;
defparam spx9_inst_4.INIT_RAM_13 = 288'h472395EF088CCAA794EAED7ABF6EAF57ABD5EAF5BEC372C160F0784CA6532983C15C2DF6;
defparam spx9_inst_4.INIT_RAM_14 = 288'h68341A0F068341A0F078341A0AF479BD5E8F37138DC8F57B411E6E37238DC2D169B91C8E;
defparam spx9_inst_4.INIT_RAM_15 = 288'h88C46253289446251178C4A6533A9D4EE774DAF5BEE171C160B0792C862EC73C8C41A0D0;
defparam spx9_inst_4.INIT_RAM_16 = 288'h2783B5BAD072C6A9D6EB5D1E40F34616C964B2697CE48655B01EB189DD3AA573C15FAB32;
defparam spx9_inst_4.INIT_RAM_17 = 288'h3854EE774BA54DE24EE662F15ABF68B49C8F68445E2D0682C1A1119954DE2B058341606F;
defparam spx9_inst_4.INIT_RAM_18 = 288'h0B7DBABB4EA858AE783C0DEE8B107DB59428E3D94C2001008080A27140E47A5E2F140D2B;
defparam spx9_inst_4.INIT_RAM_19 = 288'hDAED76BD5FB05CB0784CA6532994CA60F0571B85BEC160B0DC6E160B7D7ABD4DA6D3A9F5;
defparam spx9_inst_4.INIT_RAM_1A = 288'h371B8DE8F47A389C4E4723D1C6E371B8DC8E57A389C4D372BD9EAF583C66552B9ED3ABD5;
defparam spx9_inst_4.INIT_RAM_1B = 288'hA9D4EE9D50B960F0793CA6532590C5DD29B2A84C66310783C1A0B057AC1E11178BC1608F;
defparam spx9_inst_4.INIT_RAM_1C = 288'h44A24D28985DB39C0F38BCAA7B50B0D8AE570B6D2A71178C4A64F188C4A23118944A6553;
defparam spx9_inst_4.INIT_RAM_1D = 288'h169391EB058341A0B047A41A0F178B45206F37A40DE0EF77379A0E695D36B9599A479CA9;
defparam spx9_inst_4.INIT_RAM_1E = 288'h4883F5D4D55D95846120100C28140B09C4E27148C0F8C58D4F2994BA4C9200DE662F57EC;
defparam spx9_inst_4.INIT_RAM_1F = 288'h3C15C6C16FB0582C372B960AE370B7D7ABB4CA6D3ABF60B05BEDD5DAFD86E783C0DFAB33;
defparam spx9_inst_4.INIT_RAM_20 = 288'h168B4DC8E37138DCAF479B89C8F78C462352B9E5369B4DA6D368171B9E132B94CA653078;
defparam spx9_inst_4.INIT_RAM_21 = 288'hCBB5427B2C8E4AA31078341608F47B42231188B4160AF47ABD5EAF479B8DC8F57A389A4D;
defparam spx9_inst_4.INIT_RAM_22 = 288'hFAED2E71278BC665529944625329944A2533A9D4EA753BA6D7EC172C1E4F2794CA64B218;
defparam spx9_inst_4.INIT_RAM_23 = 288'h58240DE8F481C05FEEE6FB45ED1BA6DB2B1348F3A17AEF7FBC1E2F28245E574EAFD86C16;
defparam spx9_inst_4.INIT_RAM_24 = 288'h61389C4C261511520E895D32994A9BC4DE2DE66AFD82D37A3D1E8F58341A08F58341A0D0;
defparam spx9_inst_4.INIT_RAM_25 = 288'h0B7576994DA6D3ABD5FAFD7ABB4CA6D3EC573C1E02D94791401FCE860A2888130984C281;
defparam spx9_inst_4.INIT_RAM_26 = 288'h993C66512995CF6994B9DCC2C373C26572B95CA6530782B85BEDF60B0586E372B960AE37;
defparam spx9_inst_4.INIT_RAM_27 = 288'h58341E13188B41608F47ABD5ED057ABD5ECF579B89C2D068B49A4D372BD5E6E2723DA152;
defparam spx9_inst_4.INIT_RAM_28 = 288'hA9D4EA774BA5D329B5EAFD870593C9E4F2793C967F1564A7CB235198441A0D06834160AF;
defparam spx9_inst_4.INIT_RAM_29 = 288'hCADD1A471F7E3862D279CCE6954BA6D42C372B95C2DB4A9CCA6532994CAA553A9D4EA753;
defparam spx9_inst_4.INIT_RAM_2A = 288'h993409DECD67305A4E37A3CDE90682C0DE6F58345208F4824120903813C1DCDE68BDA354;
defparam spx9_inst_4.INIT_RAM_2B = 288'h8954F6A162B95C2DB599AC4E1EFB6BACD207D349184C260A8542815171A1670895CF2974;
defparam spx9_inst_4.INIT_RAM_2C = 288'h3C26132994CA60F0570B7DBEC161B8DC6E372B8DC6E16FAED32994DA6D369B4CA652E933;
defparam spx9_inst_4.INIT_RAM_2D = 288'h682BD5E8F57ABCDC2D068B45A8E57A3C9C6E684C6E75278C45E2F1A96D32973B9FD82E37;
defparam spx9_inst_4.INIT_RAM_2E = 288'h4C9E4F2993CFE2AC94F9E46631068341A0D068341A0B057AC223117834160AF57BC1E0F0;
defparam spx9_inst_4.INIT_RAM_2F = 288'h2B9DCAE371B756E953A9ED36B94A9D4EE7B4CA5CEE794CA5D2E994CA757EDF61B960F299;
defparam spx9_inst_4.INIT_RAM_30 = 288'h378B85C6F481BCDE9048240E06F278BB9BCD27B46675499A4460100824A6995FB0DC6E37;
defparam spx9_inst_4.INIT_RAM_31 = 288'h07EB698CA3401FCDA6C2E9BCE2834BAF9CB0995CEE953789BFDBACE60349C6F379BD20B0;
defparam spx9_inst_4.INIT_RAM_32 = 288'h1B8DC6E371B05BEBD5DA64EE793CA6D32973A9D4E24D1583C6A7D50B0DFEDB5A9BC96270;
defparam spx9_inst_4.INIT_RAM_33 = 288'h27138DCAF88D4A22D088CCA2311A9753EBF5EB7D82E372C1E0F0984C1E0AE36FB0586E57;
defparam spx9_inst_4.INIT_RAM_34 = 288'h98C42231178341E0F0683C1E11198C46233198C45E0AF47138DCCF98B3C9C2D269B91C6E;
defparam spx9_inst_4.INIT_RAM_35 = 288'hDA6D3AB74A9DCF6BB5CA65329B5FB05C70784CA68F2793CA65349A2CF62AED52A0536771;
defparam spx9_inst_4.INIT_RAM_36 = 288'h177BBDC4F6944E66F2287BC209269CD3AC796CB6572984C15FEDB4B9DCEE773DA75769B4;
defparam spx9_inst_4.INIT_RAM_37 = 288'h07F389EF299DCEA6F13783799CCF61BD1E6F47A40DE2EF6FB41A2E27241206F379BCDE2F;
defparam spx9_inst_4.INIT_RAM_38 = 288'hCA652E732994C9E29037A41E353CA6D36BB4CA5CE24B13803F9DADB6D3216EB85DB7DE30;
defparam spx9_inst_4.INIT_RAM_39 = 288'hA964FA9B5EB7D86E573C1E0F0983C15C6E161B95CAE371B0D86E160B7576994A9D4AE793;
defparam spx9_inst_4.INIT_RAM_3A = 288'h88BC1E0F068341A0D088D46A311478B45A6E371B8DC4E271B91ED068341A111994462352;
defparam spx9_inst_4.INIT_RAM_3B = 288'h1B8E0B0581C0E070584CA69347A0CE5DEC954A957A75198DCAE55288BC1A0F0995CAE552;
defparam spx9_inst_4.INIT_RAM_3C = 288'h79E54AE995CAE530781B75769B4EAF5769B4EAF57ABB4DA5D2A753A9E5329B4DAED7EC17;
defparam spx9_inst_4.INIT_RAM_3D = 288'h379385C2E279381C2E06838DE9068B4120B0481C0E02E070B8A0B189C4DE450F78C164B2;
defparam spx9_inst_4.INIT_RAM_3E = 288'h994CEE7B4CA652E73278AC0E02F07FBBDC2F382C9A492178BD60F2A9D4E24B0277B7D82D;
defparam spx9_inst_4.INIT_RAM_3F = 288'h2B95C6E572C15C6E161B0D82DF5DA5CEA752994466573CA5CEA73299445A2904824160F1;

SPX9 spx9_inst_5 (
    .DO({spx9_inst_5_dout_w[26:0],spx9_inst_5_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_5}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_5.READ_MODE = 1'b0;
defparam spx9_inst_5.WRITE_MODE = 2'b00;
defparam spx9_inst_5.BIT_WIDTH = 9;
defparam spx9_inst_5.BLK_SEL = 3'b001;
defparam spx9_inst_5.RESET_MODE = "SYNC";
defparam spx9_inst_5.INIT_RAM_00 = 288'h16934DC6E268B49A4E371BD60AF683C5E2D078CCA64F188DCB6BD60B0DCAE783C1E0F077;
defparam spx9_inst_5.INIT_RAM_01 = 288'hCBC596A953A8D3A751A8DCB255298CC6A552B954A62F1683C2A372C95CAA55298BC11C2D;
defparam spx9_inst_5.INIT_RAM_02 = 288'hEAED369D5EAED32973994CA6553CA6536BD5EB05C6E371C0E02FF7FB8DCB0794CA64F239;
defparam spx9_inst_5.INIT_RAM_03 = 288'h582C160B0481C05E2F279C162F289B48A00F282C922D2AA058F0983C1DC6FF5EAF57ABF5;
defparam spx9_inst_5.INIT_RAM_04 = 288'h68BCA251389C4DE6B22813D611299449606E068349C4E170349C9058241206F37A41A2D1;
defparam spx9_inst_5.INIT_RAM_05 = 288'hB9D4A6532894CAA773B9DCEA752A954A651268A3CDEB0583462553B9E4F277399449E4F2;
defparam spx9_inst_5.INIT_RAM_06 = 288'h89341A111993C5E0F0786D7AC161B95CF0783C1DCAE572B95CAE571B8586C572B8DFEDB4;
defparam spx9_inst_5.INIT_RAM_07 = 288'hB9DCA6331A95CAA531A8ECFE9D3D9DC9E06E067B0182D269389C2D069391E8F47B41A111;
defparam spx9_inst_5.INIT_RAM_08 = 288'hCAED7ADF60B8E06E370BFDFEDF60B8E0B0793C96433978B254A8343A9D724F0A8ECEE572;
defparam spx9_inst_5.INIT_RAM_09 = 288'h691405E7058AC5A333FA95CAE360B7D7ABD5EA757ABB4B9ED3ABD5CA5CEA7329954EE994;
defparam spx9_inst_5.INIT_RAM_0A = 288'h78AC09C2E171389C2E1723DE31278BC5E2D05834560B068AC1A2B12793C9E4F38245A4F2;
defparam spx9_inst_5.INIT_RAM_0B = 288'hB9DCEA712682C1609047A41E312A9E5369B4DA6D7ABB5EAF5729539A4D5E6500713DA312;
defparam spx9_inst_5.INIT_RAM_0C = 288'h2B9DCF0783B95CAE573B9E0AE370B0DCAE782B85B6973A9D4A6552A9D4EA732A9D4EA753;
defparam spx9_inst_5.INIT_RAM_0D = 288'h782BC9C0DF60B49A4D169345A6E683C5A0AF57C466532A964EE73288C462311EB7D82C37;
defparam spx9_inst_5.INIT_RAM_0E = 288'h0B8DCB0582C8632EF529FCBE4755B7D22372EA64EE552A954B27F41A9542BB3A8BC1A0F0;
defparam spx9_inst_5.INIT_RAM_0F = 288'hDA6D36994EAF576994DA6D36BB4CA652E973CA757ABD5FB05C2E171C0E06E17FB75BADF7;
defparam spx9_inst_5.INIT_RAM_10 = 288'h99445E2F168346251258345A24F178385E4F382C5A4B12814120B1693CAA7F50B05BABB4;
defparam spx9_inst_5.INIT_RAM_11 = 288'hCA7502C361B9DCF0782BFDAE954AABCCE00F1793DA2F1479BC9C4E479385C6F583C5E2F1;
defparam spx9_inst_5.INIT_RAM_12 = 288'h1B95CAE37FB6D32773B9DCEA773CA65264F178BC5E2F178CCA25129954EA51278BC66573;
defparam spx9_inst_5.INIT_RAM_13 = 288'h78B415ED09954AA552C9ED2E6F188D4AE6160B05C6E572B95CEE773B95CAE773C1DCAE37;
defparam spx9_inst_5.INIT_RAM_14 = 288'h1A5476635FA7D028351A8536772B954A22AF47A3DA0D0470B41A0C169345A2D57AC160D0;
defparam spx9_inst_5.INIT_RAM_15 = 288'hCA6536BD6FB05C2E170B85C70380BFDFADD6EB7D82E170B8DC6E18FC5DD6BF2C8F492AD7;
defparam spx9_inst_5.INIT_RAM_16 = 288'h280BC1C4F381C09E0F2834A2733A9E53ABF5FAF5769B4CA64F69D5EAF52E794DAF576B94;
defparam spx9_inst_5.INIT_RAM_17 = 288'h689C0E0B1482C1A08F271BCDE6F2713CDE8F78C4A6553893C62512A9D4E24F168AC52090;
defparam spx9_inst_5.INIT_RAM_18 = 288'hCA5CEA532993C5E311994CAA573A9D4EE773B9E532994DA757EC162B9E0F037FB5D26934;
defparam spx9_inst_5.INIT_RAM_19 = 288'hD9ECC6E371B95CAE572B95CAE773B9DCEE772B8DC6E572B95C6FF6EAE532973A9D4EE794;
defparam spx9_inst_5.INIT_RAM_1A = 288'h579B89C6E47ABD5E6E168341A0D168B49AD0782BD1EAF68341A152B9D4A6573CA64E2352;
defparam spx9_inst_5.INIT_RAM_1B = 288'hDAE572BB5DAF5BADF6FB85C2FD7AB2D3A570E92D9EEB63AA596C35FA7D3E814D9D49E0D0;
defparam spx9_inst_5.INIT_RAM_1C = 288'hDAFDBEBF5FAED3A9B4CA6D369B4C9DCF29B5EAED72973CA757EC170B85C2E170B85FEFD6;
defparam spx9_inst_5.INIT_RAM_1D = 288'h47AC160F1995CEA73299D4EA774BA4CE6732893C9A270178BCA050278BC5E917954EA774;
defparam spx9_inst_5.INIT_RAM_1E = 288'hDA6D369B4DA6532794CA653AA162B95C6FF6BA4CE26D279449E490482C11E6F279BC9E6F;
defparam spx9_inst_5.INIT_RAM_1F = 288'h3B9DCAE571B0D8AE572B8D82DF5EAED72973A9D4EE794B9DCEE7739944A2532A954EE794;
defparam spx9_inst_5.INIT_RAM_20 = 288'h069B9E0D0370B4DED088BC2A573994CAA553A954B27B3B995CAE572B9DCAE572B95CEE77;
defparam spx9_inst_5.INIT_RAM_21 = 288'h4A04BE6958BD6271388C2D829527834222F0783C622D0479389C4E271389C4D168B4180C;
defparam spx9_inst_5.INIT_RAM_22 = 288'hCA6D369B5CA54EA794DAF5BEDF6FBFDFEFD6DAE56E954AA5D2E974BA657ABF6FBFDF6D15;
defparam spx9_inst_5.INIT_RAM_23 = 288'hCA5D2E974893C8E04F481C0A04F281C162F299D4EE9D50B0DC2DF5EAF57A9B4CA64EE732;
defparam spx9_inst_5.INIT_RAM_24 = 288'h2B95FED74893CA6795CA449206F47A3CDE4F279BD20B078C4A2553CA54EE794DA5D2E774;
defparam spx9_inst_5.INIT_RAM_25 = 288'hFB7576994CA6536993B9DD32974A9D4A6573B9E53AA16FAED369D5DA652E732A96536A16;
defparam spx9_inst_5.INIT_RAM_26 = 288'h88BC5E311894CA22D01B95CAE783C1E0AE572B95CAE572B95C6C161B0DCAE571B0582C16;
defparam spx9_inst_5.INIT_RAM_27 = 288'h37AC1A0B047ABDA0D0579B89C2D061349A2D06730182D373415E6E372BDE0F188D4A64F1;
defparam spx9_inst_5.INIT_RAM_28 = 288'hDB656A91379BCA2753BA656E974BA6D7ADD6EB5D9A8944AC5F73FBED5616DF498B415E6F;
defparam spx9_inst_5.INIT_RAM_29 = 288'h382C5A533AA657ADF61B05BEBD5DA64EE773B9DCF29F5DA5CEE753A9D4EE994CA6536BB6;
defparam spx9_inst_5.INIT_RAM_2A = 288'h271389E8F482C1A332B9DCF2994CA6536BB5CA5D329D5BA5D2A8F2792409E70278BC5E4F;
defparam spx9_inst_5.INIT_RAM_2B = 288'hEAED36BB4DA757EC16FAED3ABF5EA5CE2512A9E5369D5FAFD7293389653EDD6A9A409E4E;
defparam spx9_inst_5.INIT_RAM_2C = 288'h3C1E0AE572B15CAE360B0582C372B95CAE571B8DC2C16FB7D7EBF60B7DBABB5EAF57ABD5;
defparam spx9_inst_5.INIT_RAM_2D = 288'h060341A0CF67B05A4E372BDA111683C2233288C46233278B4625329944560372B95CF078;
defparam spx9_inst_5.INIT_RAM_2E = 288'hA9DD36DD7DBDDE2D16AC76BF79A6BECDE0AF57B41A0D068341E0D057AC15E8F471385BEC;
defparam spx9_inst_5.INIT_RAM_2F = 288'hB9DCEE7B4FB0DBEB94A9D4EE753A9D4EA753BA6576BB5BACD1E6D26944E673399CCE6733;
defparam spx9_inst_5.INIT_RAM_30 = 288'hBA6536BB5CA6536B74B9CCD62D1589C05E0F178BC5E50382C62554DAFD82C160B7D76993;
defparam spx9_inst_5.INIT_RAM_31 = 288'hB9D4AA773CA65369D5FAF56E733EAFDBAB745893C1C0D1713CDE90584CB29B5DAE532994;
defparam spx9_inst_5.INIT_RAM_32 = 288'h3C1E0F0571B8D82C160B0582C16FB7576BB4DAFD42C361B8D82C160B0582DF5EAF57ABB4;
defparam spx9_inst_5.INIT_RAM_33 = 288'h78CCA651178C462512994CA233288AC06E572B9E0F0783C1DCAE361B0D82C15FA858AE78;
defparam spx9_inst_5.INIT_RAM_34 = 288'h679BD5ED098CC5E0D058341A08F47A3CDC6E268B45A0C060B45A2D168B45A2D57CC664F1;
defparam spx9_inst_5.INIT_RAM_35 = 288'h99CCEA774CA6532B75AA44DE4F399CCE24F27944A6775EB75FAF979B3DA2F99ED665AFD3;
defparam spx9_inst_5.INIT_RAM_36 = 288'h3803C1C0E078BC5E5058CCF29D5FB0DCAE36FAF57A9B4CA653EA371BF572973BA652E933;
defparam spx9_inst_5.INIT_RAM_37 = 288'hDAE5328F2380B81A2E1713D20F1A9E536B94BA5CEE953BA6536B74BA652A7537924162B1;
defparam spx9_inst_5.INIT_RAM_38 = 288'hEAED769B4EAFD86E371B8DC6E370B0582C160B7DBEBD5CA5CEE752B9ED36BD5EAE52A7D5;
defparam spx9_inst_5.INIT_RAM_39 = 288'h580DC6E572B9E0F0783B95C6C360B057EBF51B15CF0984CA64F0571B8DC6E370B05BEBD5;
defparam spx9_inst_5.INIT_RAM_3A = 288'h270B45A2D169345A2D269349C4D168B49CD088C45E31188BC6651158342A573B9C4622F1;
defparam spx9_inst_5.INIT_RAM_3B = 288'h99CCE6954BA6DBF0390CE5D68333A4DFB5DA8BF4D5E8F57B41E13188B411E8F479B89C4E;
defparam spx9_inst_5.INIT_RAM_3C = 288'h2B9DC6FF6FA85BEBB5DA7D42DF5DA6D369B4DADD26733A9D52E974AA552E9549A4D2A954;
defparam spx9_inst_5.INIT_RAM_3D = 288'hB9DD2A733A9D4EA753A9DD2E953AA4CE66F248240E070380BFDDEE178BC9EB1A9F57ADD5;
defparam spx9_inst_5.INIT_RAM_3E = 288'h0B0DCAE371B0D82DB4B9DCE6553CA6D369B4CA6532953A9DD264D1378B89C2E27AC2A773;
defparam spx9_inst_5.INIT_RAM_3F = 288'hFAFD7EA362B9E132B95CA60F0582B8DC6E160B7DBABD5EAF57ABB5EAFDBEC160B0582DF6;

SPX9 spx9_inst_6 (
    .DO({spx9_inst_6_dout_w[26:0],spx9_inst_6_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_6}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_6.READ_MODE = 1'b0;
defparam spx9_inst_6.WRITE_MODE = 2'b00;
defparam spx9_inst_6.BIT_WIDTH = 9;
defparam spx9_inst_6.BLK_SEL = 3'b001;
defparam spx9_inst_6.RESET_MODE = "SYNC";
defparam spx9_inst_6.INIT_RAM_00 = 288'h2723DA0F0683C1E2D078C45E2D078D4F69B4CA4CA23110B0D86E572B9DCF0783B9586C15;
defparam spx9_inst_6.INIT_RAM_01 = 288'hFD7EA2FD3579B9E151A9445A0D0683411E4D068345A2D06834180D068345A4D269345A2D;
defparam spx9_inst_6.INIT_RAM_02 = 288'hEAF57AB94AA54EA753BA5D2673399D52A975BAD52A9139A65830390C75F2D35598482537;
defparam spx9_inst_6.INIT_RAM_03 = 288'hAA4496290481C162F23803B9DCEF70BD6333CAF57ABF5FAFD7EBF5EAED32973CA6D369F5;
defparam spx9_inst_6.INIT_RAM_04 = 288'hDA7D7ABD5DA54E653299CCDA24F170B89E6F68CCEE753A9D4EE97499C4E673399CCEA774;
defparam spx9_inst_6.INIT_RAM_05 = 288'h2C15C6E16FB7D7ABD5FB0582E371B95C6E170B7D82C160B0D82DF6FAF572993DA6D369B4;
defparam spx9_inst_6.INIT_RAM_06 = 288'hB9E5329539944663D5FB0586E572B9E130783B9582BF5FAFD42C573C26132B94CA653078;
defparam spx9_inst_6.INIT_RAM_07 = 288'h579B85A0D060341A0C06834180C060B49A4D168341A6E7844622F1582BD60F178B41A0F1;
defparam spx9_inst_6.INIT_RAM_08 = 288'hAAE576D96BAEDBEFF7EBEDB6FB6AABD0E4525A55F33DADCA56A28F57C4262F047A3D5ED0;
defparam spx9_inst_6.INIT_RAM_09 = 288'h071C1E574EAF57ABF5EAF576993B9D4EE793DA757ABB5DAF57295399D52E974BA5526954;
defparam spx9_inst_6.INIT_RAM_0A = 288'h27A41A2F18954EA753A9DD3295399C4A2533A9DD2E97489345A2B138241A49027FBB5BAD;
defparam spx9_inst_6.INIT_RAM_0B = 288'h1B8DC6E572B95CAE571B7DBEBF5EAED369B4DA6D369D5FAFDBEDF5EADCE24F2792C0DE4F;
defparam spx9_inst_6.INIT_RAM_0C = 288'h2B9DCF0773B8D86C160B0D86E573C26132B95CA64F0782B8DC2C160B0DC6E371B8DC6E37;
defparam spx9_inst_6.INIT_RAM_0D = 288'h169349C2DF6034DCF198C4622D047AC222D068345A111994CA231188CCB6BD5FB0D86E57;
defparam spx9_inst_6.INIT_RAM_0E = 288'h49A4DEB78ECE66B117F9BBD1CAF783411E6E47ABD5E6E371385A0D06833D82D067B3D80C;
defparam spx9_inst_6.INIT_RAM_0F = 288'hA954F27B4DAE5329B4DAD4E6733AA552A955BAD56AB55CB7DFF1F7FB863F1B7BACD1E6B3;
defparam spx9_inst_6.INIT_RAM_10 = 288'h8944AA753AA5D2A73399CCDE4B1382C5227007EB6D9AC17B46E9D5EAF57EBF5EAE52E753;
defparam spx9_inst_6.INIT_RAM_11 = 288'hDAED36994DA6D3ABD5FA8582C16CA449E2D1581BC9E4F5844A24F19954EA753BA652E933;
defparam spx9_inst_6.INIT_RAM_12 = 288'h3C26130994C1E0F0782B8DC6E573C1E0F0582C15C6E371B95CAE573C1E0AE370B0582DD5;
defparam spx9_inst_6.INIT_RAM_13 = 288'h684C5E2F178ABD5EB068445E2F1A96D7ABF60B0D86E572B9DCF0772B95CAE361B0DCAE78;
defparam spx9_inst_6.INIT_RAM_14 = 288'h57ABD5EAF479389C4E271381A0C060305A0CF67B3D82D271B85A2D271B9A0D068445E2D0;
defparam spx9_inst_6.INIT_RAM_15 = 288'h89C4E69559AD56AB96FC0E473B7BADD72D969AB4D26B49B66373388BBD8A930168B51EAF;
defparam spx9_inst_6.INIT_RAM_16 = 288'h48A44E00FD6D2E97CD68DD36BB5DAFD7EBD5EA64EE773B9E4F2994CA65329748944E6713;
defparam spx9_inst_6.INIT_RAM_17 = 288'hA9BC560903793C5C9079449E312A9CCEE994BA5D2A73399CCE6753BA4CEA974BA55224B1;
defparam spx9_inst_6.INIT_RAM_18 = 288'h3C1E0F0983C0DC2C371B8D82C161B0D86E371B8DBAB94DA6D369B4DA64EE7D50B7D7AB94;
defparam spx9_inst_6.INIT_RAM_19 = 288'hEAF57EC160B0586C572B9DCEE773B95CAE361B95CAE783C1E0F0783C26532782C15CB078;
defparam spx9_inst_6.INIT_RAM_1A = 288'h06033D80C067B05A4D2723DA0D057ABD5EB0682BDA0F178C46231188BC5E2F188C45E311;
defparam spx9_inst_6.INIT_RAM_1B = 288'hCB6DF2F56BB6E370F6198CCA85409EC95E0D169B95ECF57A3D1E6E271B89C2D06830180C;
defparam spx9_inst_6.INIT_RAM_1C = 288'hEAF5769D5DA6D32993B9DCF2994BA4CDE4D27944E26F369B4DA6F3BB7E3F176AADDB2D96;
defparam spx9_inst_6.INIT_RAM_1D = 288'hB9E532974A9D4EA753895532B94AA5D2E954BA44D229158943DDADA6533DCD1A9DD2E794;
defparam spx9_inst_6.INIT_RAM_1E = 288'h0B0586E571B85BEBF5FAF5727318844729F5EAE52A733892C09E0E0703920F278C4A2533;
defparam spx9_inst_6.INIT_RAM_1F = 288'h3B95C6C161B15CAE572B95CB0784C260F0783C1E0AE371B95CAE37FB7D7EBF60B0582C16;
defparam spx9_inst_6.INIT_RAM_20 = 288'h47A3D60D0583C222D078C46233288BC6231188CCA6594DAF57EBF5FB0586C372B9DCF078;
defparam spx9_inst_6.INIT_RAM_21 = 288'hB8BBD1C6E271B8DC6E3723D1E6E370B7D9ECF60341A0C060B45A0CF67B05A6E57BC1E0D0;
defparam spx9_inst_6.INIT_RAM_22 = 288'h89349A4D269349249269D5AED769ACD62955CB6DF6F96BB65F71979B3542791B8ECBE7D2;
defparam spx9_inst_6.INIT_RAM_23 = 288'hCADD2A974792456291287BAD96CD68BDA353BA65369D5DA6D369B4DA652E753A9DD2A733;
defparam spx9_inst_6.INIT_RAM_24 = 288'h995CF6994CA652A712580BB59CD17241A2D18944A6794BA54E6753A9DD2E974CAE572B95;
defparam spx9_inst_6.INIT_RAM_25 = 288'h3C160F0783C160AE371B8DC2DF6FAFDBEC161B85BEBF61B0DC6E360B7576993A9445E111;
defparam spx9_inst_6.INIT_RAM_26 = 288'h78C45E311994CAA774DAF57ABF50B0586C573B9E0F0783B95C6C361B8D82C361B95CF078;
defparam spx9_inst_6.INIT_RAM_27 = 288'h16FB3D80C06030180C168B419ECE5830DCAF68341A0AF58341A0B0683C5A0F188CCA6511;
defparam spx9_inst_6.INIT_RAM_28 = 288'h493CE6B55BB6DF6F96BBD5E2C7409F4B6391D974B65307833D1E4E068B49C6E47A3D1E6E;
defparam spx9_inst_6.INIT_RAM_29 = 288'h27AC66573CA7576BB4CA6D3ABB4CA54E6753A9CCE26F2692C52291593CE2935BB65A6AB2;
defparam spx9_inst_6.INIT_RAM_2A = 288'h382C5A3129954F2974A9D4EE974BA6576B95CAE576B95BA552E8F358AC52250E75331BEE;
defparam spx9_inst_6.INIT_RAM_2B = 288'hFB7D82C360B7D42C571B0582C16EAE4EA4F0784CAE773CA65369D5EADCDE290076B3582E;
defparam spx9_inst_6.INIT_RAM_2C = 288'h0B0DCEE784C26130783B95CAE361B0582C160B0DC6E571B8DCAE572B95C6E370B7D7ABF5;
defparam spx9_inst_6.INIT_RAM_2D = 288'h060B4DCAF579B91EF188BC11EAF68342655299446231178C45E2F0783CA6774CA6D7EA16;
defparam spx9_inst_6.INIT_RAM_2E = 288'h2A74B63F2C8BBD1C8E371389C2D169389C6E271389C2D067B019ECF67B0180C168B419EC;
defparam spx9_inst_6.INIT_RAM_2F = 288'h894CE67339A4CDE491489C52514DBF632CD359B4DE8D359249A534DB86433773984928B5;
defparam spx9_inst_6.INIT_RAM_30 = 288'hBA6572B95CAED72B74AA55266D2489C41FAED6EB7DC7058BCA6774DAED72994DAFD7AB74;
defparam spx9_inst_6.INIT_RAM_31 = 288'hDA64F2994DA6D329B4EAFD7EDD5B9BC5200EE6F37DA2F58C4A2533AA5D32994CAED6E954;
defparam spx9_inst_6.INIT_RAM_32 = 288'hFAF57ABD5EAFDBEDF6FB0582C160B7DBEDD5DAE536BD5FA8582C361B0DC6C16FB0586DF6;
defparam spx9_inst_6.INIT_RAM_33 = 288'h784CAA73268341A0F1B9DCEE793583C66774DA757EC162B95CF0984C26130983C15C6E16;
defparam spx9_inst_6.INIT_RAM_34 = 288'h271385A0DF67B09C6E268B7D7CBF6033D9EC060B49A4D3723D1E4E16939E13178C466511;
defparam spx9_inst_6.INIT_RAM_35 = 288'hAB65A6AD328FBFDE3079EDC7219CBD5AEF164A04CA813E97CBA50F160301A2D169389C4E;
defparam spx9_inst_6.INIT_RAM_36 = 288'h287BF5D8DE70C162D1895D32994CA6532994EAE526733BA55266F3692C4E2918A65B2F35;
defparam spx9_inst_6.INIT_RAM_37 = 288'h892401DADD66B45EB18944E6753CA656E974BA4CE6774BA5D2E954BA552A974BA4D1A491;
defparam spx9_inst_6.INIT_RAM_38 = 288'hFAFDBEDD5EAF57EC160B0586C361B0D82DF6EAF57ABF5FAFD7ABD5FAF5769D5EAED72953;
defparam spx9_inst_6.INIT_RAM_39 = 288'h68C4AA794DAF57EC161B95CEE784C26130983C15C2DD5DA65329B5EAFD7EBF60B05BEDD5;
defparam spx9_inst_6.INIT_RAM_3A = 288'h067B0184D271B8DC8E57A385A0D37B41E0F0995CEA51188CCA64F178B41E352994CA646F;
defparam spx9_inst_6.INIT_RAM_3B = 288'hBBC5528530984FE7D2C8C3C99EBF67B05A4E27134DC8E3703799CBE5934DC4D16833D9EC;
defparam spx9_inst_6.INIT_RAM_3C = 288'hCA5CEE994BA44A2554AA4CE26F389CD2EB76CB6DE6AD3491479F4DC6ACAEDD8FC7E7B197;
defparam spx9_inst_6.INIT_RAM_3D = 288'hBA54E6733894CEE974AA552A933AA5D32B95AA3CD6230D76375DEF38349A512A9E532994;
defparam spx9_inst_6.INIT_RAM_3E = 288'h0B0582C16FAFDBEDF5EAF57ABD5EAF57ABB4BA5CEA7326893FDB8CC67B4E0F299DD32994;
defparam spx9_inst_6.INIT_RAM_3F = 288'h3B9DD30983C0DBEBD5DA6D369B5EAF57ABF5FAF57ABD5FB0582C160B0DC6E371B8DC2C16;

SPX9 spx9_inst_7 (
    .DO({spx9_inst_7_dout_w[26:0],spx9_inst_7_dout[8:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_7}),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[8:0]})
);

defparam spx9_inst_7.READ_MODE = 1'b0;
defparam spx9_inst_7.WRITE_MODE = 2'b00;
defparam spx9_inst_7.BIT_WIDTH = 9;
defparam spx9_inst_7.BLK_SEL = 3'b001;
defparam spx9_inst_7.RESET_MODE = "SYNC";
defparam spx9_inst_7.INIT_RAM_00 = 288'h57A3D5F119954AA51188CCA2332993C5E2D05823D62D168C4AA794DAF57EC161B15CAE57;
defparam spx9_inst_7.INIT_RAM_01 = 288'h06934DC4D269B8DC6E0672F97EC060B41A0D168B419EC060B4DC8E479B8DC8F371389CAF;
defparam spx9_inst_7.INIT_RAM_02 = 288'hBAEDEED358A2CFE10C75DB420D3DB96875B8BBDDEEF364A048245419FCF22AD05F2BD60C;
defparam spx9_inst_7.INIT_RAM_03 = 288'hCAE572B5489AC81F8DB6EB7DC5058B49E533BA6D7ABB5CA5D2E9338944A6754AA5D2A955;
defparam spx9_inst_7.INIT_RAM_04 = 288'hFAF572973B9DCE64F25803B198CD68396333CA656E97499BCA271289CCEA933AA5526774;
defparam spx9_inst_7.INIT_RAM_05 = 288'hDAF57ABF6FB7DBEDF6FB0582C161B0D86E572B8DC2C361B0DC6E160B7D7ABB4DA65329D5;
defparam spx9_inst_7.INIT_RAM_06 = 288'h78B4160B06824562D1894CAA794DAF542C161B0D86C362B9DCF0782B8582BF5EAED369B4;
defparam spx9_inst_7.INIT_RAM_07 = 288'hE5FB0182D16FB3D80C169B95ED0479389C6E57ABD60AF37938DED09964EE532993C6E773;
defparam spx9_inst_7.INIT_RAM_08 = 288'hDC65F2F778A9CC22744A9D06654C8AB7D5EBF58305A2D268B45A6E270341BECF67B3D9CC;
defparam spx9_inst_7.INIT_RAM_09 = 288'h793CA67B5FB05C2DF6CACCDA4D1AA5D32B95BADD668B27A4D5A9CF963AE9BF08AF6075F9;
defparam spx9_inst_7.INIT_RAM_0A = 288'h17AC62553BA5D2E953793CA26F258CCEA954AA5D2EB75BAE56A91348FBF1B4CA66B41E91;
defparam spx9_inst_7.INIT_RAM_0B = 288'hFB0582C372B95C6E371B85BEBD5DA6D36993B9DCF69F5EAED36994BA54DE4B027F3719AD;
defparam spx9_inst_7.INIT_RAM_0C = 288'hDAFD42C361B0D86C361B0D8AE571B0D82DF5EAED7ABF60B05C6E371B85C2DF6FB05BEDF6;
defparam spx9_inst_7.INIT_RAM_0D = 288'h169385C6E683C15E6F47938DEF0A94CA6552A95CE22AF684CAA552E6A46275499D4EE994;
defparam spx9_inst_7.INIT_RAM_0E = 288'hF57289A2D067B05A6E47238DC4D06833D9ECF603019ECE5F2FD9ECF6034DCAF67ABD5E6E;
defparam spx9_inst_7.INIT_RAM_0F = 288'hBA5D266B279CD6AAB3085BA9A308AEE3F219EC65EEF779B253E3D0091D128D54AFCA5E8D;
defparam spx9_inst_7.INIT_RAM_10 = 288'h89D52A933AA4CE6974BADD266D2F7DB6D94CF79C5A51389D536BD6EAED6E933692412333;
defparam spx9_inst_7.INIT_RAM_11 = 288'hEA6D3A9D5EAF57ABD5EAED7ABD5CA54DE4B127EB297ED6944E673399DD2A8F27944DE4D2;
defparam spx9_inst_7.INIT_RAM_12 = 288'h1B0DC6C361B8DC6E571B8DC2DF6FB7DBEDF6FB7DBEBD5EAFD42C160B7DBEDF5EAF57ABD5;
defparam spx9_inst_7.INIT_RAM_13 = 288'h88CCAA55288B411ED0A964EE470694D32BF7FBFDFEDF6FB0586C362B1586C360B0582A16;
defparam spx9_inst_7.INIT_RAM_14 = 288'h168B419ECF603019EBE5F2F980D3723D5EAF47ABD1E2D3723D60F0682BD1EAF47A3DA111;
defparam spx9_inst_7.INIT_RAM_15 = 288'h2D06771779B350E611D853F60736AA5067B17702F55AAF59B4DA2D062395EAF471341A0D;
defparam spx9_inst_7.INIT_RAM_16 = 288'hD773B5C0F5944E2733BA6532974A9C4DE4914834A6754AA4D269158A350A25159D5BF05A;
defparam spx9_inst_7.INIT_RAM_17 = 288'hA9D4E66B1E6D2FDAB17944E6754BA552671379349E513AA552693389C4EEB75BA4D1A5EE;
defparam spx9_inst_7.INIT_RAM_18 = 288'hEAFDBEDD5EAF576BD5EAFD7EBF5FB7DBABB4DA6D369B4DA757EBF5FB7DBEBD5DAED76974;
defparam spx9_inst_7.INIT_RAM_19 = 288'h6944B2BD60B960F2994C9E130984C1DC6C360A8542C362B95CAE572B960AE37FB6D76BB5;
defparam spx9_inst_7.INIT_RAM_1A = 288'h471385A6E57A3C9C8F58341A08F47ABD60B068341A0F188C45E2D0683C1A111A94C8E291;
defparam spx9_inst_7.INIT_RAM_1B = 288'hE93B817A9D4EAB960C472391C6E57ABCDC2D067B3D82D16837D9EC06033D9CBE5FB05A8E;
defparam spx9_inst_7.INIT_RAM_1C = 288'h89BC962B189D52A9349A6DEECF44934F2E3A5E26CB5D8AB351A8B408D3A5DD0199D0E854;
defparam spx9_inst_7.INIT_RAM_1D = 288'hBA55266D2593CA2754AA552A9339A5D6EB559A348600F07FBC60B289CD2A974BA552A733;
defparam spx9_inst_7.INIT_RAM_1E = 288'h0B7DBABB4DA6D32994EA757ABF60B7D7ABB4CA5D2E753A9D4DE40ED683920B1794CEE974;
defparam spx9_inst_7.INIT_RAM_1F = 288'h5CA60EE573B95CF0783C1E0B0582B8DC2DD6DAE532994CA65329B4CA6D36BD5EAF57EC16;
defparam spx9_inst_7.INIT_RAM_20 = 288'h57B41A0F0682BDA0D068341E332B94C5E0F0988385E6F483CAE9F63C2E9F6FB6D369B4B9;
defparam spx9_inst_7.INIT_RAM_21 = 288'h26FB397CCE6733D80C068345BECE5F2C182D168B45A4E168349C6E37A3C9C2E2723CDC8F;
defparam spx9_inst_7.INIT_RAM_22 = 288'h2D1ECF65BDC455EB1539EBE1B8FF894D6AD53A6C59C2BD56A795EBF58309AAE77BBD5E8E;
defparam spx9_inst_7.INIT_RAM_23 = 288'hBAE56A93489AC861EFE78C0E2F3BAD52A974BA5D2E95499BCA2754AA4CE2714AAD572DF8;
defparam spx9_inst_7.INIT_RAM_24 = 288'hDA6D369B4DA652A75399CCD200E17A4162D289552E974AA4CDE4D2794D2A93399D52A954;
defparam spx9_inst_7.INIT_RAM_25 = 288'h1B85BEDD5CA5D2A733994CAE794DAF576BB5FA8582DF6EAED7ABD5EAED2E794DA6D3A9B4;
defparam spx9_inst_7.INIT_RAM_26 = 288'hA954AA351C60392133BA6D7EC162BA6574DA6D2E972BA6D369B4DA6D36974B94CA64F058;
defparam spx9_inst_7.INIT_RAM_27 = 288'hE58B4DC4E168345A2D168B49C8F47ABD1E6E47ABDA0F057B41A0B0682C15EAF57B422331;
defparam spx9_inst_7.INIT_RAM_28 = 288'h3A7CB210F46FAF1369E51315D10883BD5C8E268B0180CF6733D9ECF67B399CC060B7D9AB;
defparam spx9_inst_7.INIT_RAM_29 = 288'hBADD2E954A9CCE675499D4EA91389D536DF70C0E4B25A0CEE2EF776A7C71FD0292D1AAD5;
defparam spx9_inst_7.INIT_RAM_2A = 288'h482C5A513AA5D6A9339A4CE271389CCE69349A5D72B95CADD668F3388C06030080C1A575;
defparam spx9_inst_7.INIT_RAM_2B = 288'hEAED76BD5FB05BEDD5EAF57ABD5C9D4AA573B9ED36994CA65369B5CA5CEA774CAD51220F;
defparam spx9_inst_7.INIT_RAM_2C = 288'h3C26532B95D369B4BA5CA6130783C26172B94CA64F037FB5D2A71278C4AA794DAF5BEDF6;
defparam spx9_inst_7.INIT_RAM_2D = 288'h57A3D1EAF683C1E2D057ABD5EB0379B91E6E57BC22332A954AE56BF69BDE353DA7D86E57;
defparam spx9_inst_7.INIT_RAM_2E = 288'h5713419ECF672FD9ECF6030180CF672F97ECF67B397CB168B45A0D068B49C2D06938DC8F;
defparam spx9_inst_7.INIT_RAM_2F = 288'hEB0E0725A2D067F1B89B2CD2631E86C064944A14FE5705682F940B362355CCE77BBE20F0;
defparam spx9_inst_7.INIT_RAM_30 = 288'h9A5526934BAE572B75AA44D64301814061CEF7ACB2BB5CADD2A93399CCEA933793C9E754;
defparam spx9_inst_7.INIT_RAM_31 = 288'h994CA6552B9DCEE773CA6532994BA5D32BB5DABC85E9148AC9E533AA55269549A4CE2713;
defparam spx9_inst_7.INIT_RAM_32 = 288'h3B9E0F0582B95C6E17FB7572953893CA6753BA6D7ADF60B8DC2E16EAF57ABF5EAF576B73;
defparam spx9_inst_7.INIT_RAM_33 = 288'h379B89C8F783C5E0F098DC7980D272C26574EAFD82C372B95CB0784C26572B95CA64F077;
defparam spx9_inst_7.INIT_RAM_34 = 288'hF67B397CCF67B3D9ECF67B3D80D271385A0D271B8DC6E371B95E8F57BC222AF47AC11E6F;
defparam spx9_inst_7.INIT_RAM_35 = 288'h2914FA30F260AC986C361311AEE87CC2610F4713419ECE5FAFD80CE5F2F97EC0603019EC;
defparam spx9_inst_7.INIT_RAM_36 = 288'h087BEDBCE6975BAD95BA552A95399D51E49158C4F2A182C8E47219EC6DF2F36194B5D98F;
defparam spx9_inst_7.INIT_RAM_37 = 288'hCAED72BB5899C1209158B4A2734BADD6A93389C4E2754AA4D2EB54AA55226D2591C41FEF;
defparam spx9_inst_7.INIT_RAM_38 = 288'h99BC5A2D1795536C171B8DC2FD6EB7DBABB5DAED32953994CA65328944A6574CA5D2E794;
defparam spx9_inst_7.INIT_RAM_39 = 288'h58446A593DA753ABF50A8582C161BA6174DA6D36972983C15C6E361B8DCB0793C0E3ED94;
defparam spx9_inst_7.INIT_RAM_3A = 288'h067B0184D371B89A6E47ABC9C4E685495E8F68341E0D057A3CDCD098ABDE111880B45C6E;
defparam spx9_inst_7.INIT_RAM_3B = 288'h160B0580CF67B019ECE5F2FD7CBE5FB0180C060B45A2D06733962D26837D80C067B01A0D;
defparam spx9_inst_7.INIT_RAM_3C = 288'h792C964F3AA6D830390C6DF6FF8EC65E2BF1760A4124B36130562C77542E17097B391A4D;
defparam spx9_inst_7.INIT_RAM_3D = 288'hCB5D627139A4D2691389DD6A93389AC461CEC6D331BAED74301F34FBFDF6D75AA552A953;
defparam spx9_inst_7.INIT_RAM_3E = 288'h1C756E773BA5CEE753A9CC9E2B05844AA773CA6536BD6FB75B2B133814122B27944EA995;
defparam spx9_inst_7.INIT_RAM_3F = 288'h0B0D8AE786D3EDF6DA5CA60F0782C160B0370B85C70591C75AA8B138241A333CA8DD3299;

SP sp_inst_8 (
    .DO({sp_inst_8_dout_w[30:0],sp_inst_8_dout[9]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9]})
);

defparam sp_inst_8.READ_MODE = 1'b0;
defparam sp_inst_8.WRITE_MODE = 2'b00;
defparam sp_inst_8.BIT_WIDTH = 1;
defparam sp_inst_8.BLK_SEL = 3'b000;
defparam sp_inst_8.RESET_MODE = "SYNC";
defparam sp_inst_8.INIT_RAM_00 = 256'hFC0007000000000000003003E3FFFFFFFFFFFFE00000FC783FFF0020F0000000;
defparam sp_inst_8.INIT_RAM_01 = 256'hBC000780003FFF90207000000000000003003EFFFFFFFFFFFFFC00003F8E03FF;
defparam sp_inst_8.INIT_RAM_02 = 256'hFFFFFE7FFFFFFF9800000303FFFF0F07800000000000003007FFFFFFF7FFFFFF;
defparam sp_inst_8.INIT_RAM_03 = 256'h00000000001BFFFFFFFFFFFFFFF70001FFF87FFFF0F0380000000000000000FF;
defparam sp_inst_8.INIT_RAM_04 = 256'hFFF8463C0000000000000103FFFFFFFFFFFFFFFFC000FFFF1FFFFF8F03C00000;
defparam sp_inst_8.INIT_RAM_05 = 256'hFF300FFFFE1FFFFF80F3C000000000000018DFFFFFFFFFFFFFFFF8003FFFE3FF;
defparam sp_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFDFE03FFFFE3FFFFF81F9E000000000000019FFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_07 = 256'h0000000003FFFFFFFFFFFFFDFC7FC07FFFFE3FFF9FC000F00000000000001FFF;
defparam sp_inst_8.INIT_RAM_08 = 256'hFFFFE0F07C0006000000003FCFFFFFFFFFFFA7CFF01FFFFFC3FFFFFC06078000;
defparam sp_inst_8.INIT_RAM_09 = 256'h3FF83FFFFE07FFFF9F9FC0E001800000000FF9FFC7FFEFFFF031FFC1FFFFF03F;
defparam sp_inst_8.INIT_RAM_0A = 256'hFF0F1E1FFC0001FF07FFFFC07FFFE3F1780E018004000003FF3FF878F8FFFC02;
defparam sp_inst_8.INIT_RAM_0B = 256'h000000019FFE7FE0C1CFFF80003FE07FFFFC0FFFFFFF0780F02007C000047FEF;
defparam sp_inst_8.INIT_RAM_0C = 256'hFF9FFFE1FC78000000003FFFCFFC0039FFF00003FC07FFFFE1FFF3FFFF07E780;
defparam sp_inst_8.INIT_RAM_0D = 256'h07E019BFFFC3FFF9FFFE7FFF81C0000007FFF0FF80077FFE00003F80FFFFFC1F;
defparam sp_inst_8.INIT_RAM_0E = 256'hFE001BFFF80000F8007FFFF83FFFCFFFC1FDFC700600007FFE9FF000FFFFC000;
defparam sp_inst_8.INIT_RAM_0F = 256'hC01FF0001FFFFFC0027FFF80001E00FF9FFF03FFFCFFF33FFF9E01F00003FFFF;
defparam sp_inst_8.INIT_RAM_10 = 256'hFFFF3F1FFFFFFDE1FF0003FFFFC8000FFFF00001C01FF3FFE07FFFFFFC7FFF7F;
defparam sp_inst_8.INIT_RAM_11 = 256'h07FFFC07FFE1FFFFFFFFFE7FBF7C1FE0003FFFF80003FFFE00003E03F83FFF0F;
defparam sp_inst_8.INIT_RAM_12 = 256'hE0030FFFE00000FFFC007FFC7FFFFFC7FFE1FFDFC0000007FC3F00083FFF8000;
defparam sp_inst_8.INIT_RAM_13 = 256'hFF0000E007E01C0061FFF800001FFE0007FF8FFFFFF87FFF1FFFF80000407F03;
defparam sp_inst_8.INIT_RAM_14 = 256'hFFFFFF7FFE1FFE01000E00F80080047FFA100000FF00007FF1FFFFFFF7FFE1FF;
defparam sp_inst_8.INIT_RAM_15 = 256'h03C00007FF87FFFFFFF9FC387FC00000E03F000000DFFF4000001F80000FFE3F;
defparam sp_inst_8.INIT_RAM_16 = 256'h00011FF80000F060007BC3F8FFFFFFFF9F83CFF800000C7FF0000019FFC80003;
defparam sp_inst_8.INIT_RAM_17 = 256'h0003C3C3FFC0000023FF0019FC000F9FF8FF9FFFFFFE787EFDF80000001FFE00;
defparam sp_inst_8.INIT_RAM_18 = 256'hFFFFFFFE7FF807FFF9FEFFF80000003FE007FF803FE3F807F3FFFFFFEFE7FFC0;
defparam sp_inst_8.INIT_RAM_19 = 256'h0F811F803F87FFFFFFF7F1FF07FFFFFFFFFF00000004FD80FFF01F0CFE007C7F;
defparam sp_inst_8.INIT_RAM_1A = 256'h000003F807FF8FC047E007F9FFFFFFFFFF1FE0FFFFFFFFFFF00000001F701FFC;
defparam sp_inst_8.INIT_RAM_1B = 256'hFFFC0001FFC00700007E01FFF3E019F800FF3FFFFFFFFFFBFC1FFFE000FFFE00;
defparam sp_inst_8.INIT_RAM_1C = 256'hFFFFFFFFFE73FFFF00001FF800F00007003FBFE0027E001FE7FFFFFFFFDFFF9F;
defparam sp_inst_8.INIT_RAM_1D = 256'h0033E0007F9FFFFFFFFFFFF0FFFF80000006000F0000C007E3F000CF0003FCFF;
defparam sp_inst_8.INIT_RAM_1E = 256'h078000003C07000C78000FE3FFFFFFFFFFFF0FFFF8000000000078000001F03C;
defparam sp_inst_8.INIT_RAM_1F = 256'hFFF00F03F800003C00000780C0031E0001F87FFFFFFFFFFFF3FFFF8060000000;
defparam sp_inst_8.INIT_RAM_20 = 256'hFFFFFBFFFFFFFFFE0078FFFE0007E00000F010008780003C1FFFFFFFBFFF9FFF;
defparam sp_inst_8.INIT_RAM_21 = 256'h387000007E7FFFFFFFFFFFFCFFFFE007CC1FFF007C00001E020061E00001E3FF;
defparam sp_inst_8.INIT_RAM_22 = 256'h00F8000030081C1C00001FCFFFFFFFFFFFFF9FFEFC003CE007F0078000018040;
defparam sp_inst_8.INIT_RAM_23 = 256'hF7F80C3C3800300F00000E03FE0F80000FF9FFFFFFFFFFFFF7FFDF8087C70003;
defparam sp_inst_8.INIT_RAM_24 = 256'hFFFFFFFFFFFFFCFF8001E1C00200E00001C07C03000001FF1FFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_25 = 256'hF800000FF8FFFFFFFFFFFFFBFF9FF0001E1F00201C0000180C03E000003FC7FF;
defparam sp_inst_8.INIT_RAM_26 = 256'h40380C006041FC000007FF83FFFFFFFFFFFF3FF7FC0000C07C1E038000030007;
defparam sp_inst_8.INIT_RAM_27 = 256'hFFE0000000060006000000083F800001FFF83FFFFFFFFFFFE3FFFF80000003FE;
defparam sp_inst_8.INIT_RAM_28 = 256'hFFFFBFFFFF9FFFFC0000000000000000000007E000007E7F03FFFFFFFFFFFCFF;
defparam sp_inst_8.INIT_RAM_29 = 256'h000007F0FC67FF1FF7FFFFF3FFFFC0000000000000000000007800000F8FE03F;
defparam sp_inst_8.INIT_RAM_2A = 256'h000000000000000007F83F1C6C3FFFFFFFFFFFFFF00000003F8000000000000C;
defparam sp_inst_8.INIT_RAM_2B = 256'hFFE00000001E000000000000000001FC006380EFFFFFFFFFFFFFFE00000001F0;
defparam sp_inst_8.INIT_RAM_2C = 256'hFFFFBFFFFFFFFFFF00001001C000000000000E0000000000201FFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_2D = 256'h040000000007FFFEF3FFFFFFFFFFF080010000000000000000C000000000001F;
defparam sp_inst_8.INIT_RAM_2E = 256'h000000000007018000000001FFFFFFFFFFFFFFF7FFF03FE00000000000000038;
defparam sp_inst_8.INIT_RAM_2F = 256'h1FFF801EFE00000000000300E420000001807FFFFFFFFFFFFFFCFFFC03FF8000;
defparam sp_inst_8.INIT_RAM_30 = 256'hFFFFFFFFFE7FE3FFF07FBE000000000000380000000003801FFFFFFFFFFFFFFF;
defparam sp_inst_8.INIT_RAM_31 = 256'h0000004000FFFFD9F7FFFFC7FFFFFFFFFF8000000000000700000000000003FF;
defparam sp_inst_8.INIT_RAM_32 = 256'h000000000F0000000060001FFFFF1FFFFFF8FFFFFFFFFFFE0070000000007000;
defparam sp_inst_8.INIT_RAM_33 = 256'hFFFFFF0FFC000000000003E0000000000007FFFFDBFFFFFF1FFFFFFFFFFFC008;
defparam sp_inst_8.INIT_RAM_34 = 256'h9FE7FFFFFC0FFFFFFFE1CF8000300000007800000000001FFFFC7F3FFFFFE07F;
defparam sp_inst_8.INIT_RAM_35 = 256'h000000607FFFFA3EFFFFFF81FFFFFFF83BF000060000000F000000000007FFFF;
defparam sp_inst_8.INIT_RAM_36 = 256'h1C0000007800000006300FFFF3C4FFFFFFF01FFF007807F60000E0000001E000;
defparam sp_inst_8.INIT_RAM_37 = 256'hFC0007FFF00003C000000F000000038003E3FC7CBFFFFFFE01FFE00C01FE0000;
defparam sp_inst_8.INIT_RAM_38 = 256'h39FFFFFFF803FFE0007FFF800038000001E0000003C60079FF8FEFFFFFFFC01F;
defparam sp_inst_8.INIT_RAM_39 = 256'h006103073BFC607FFFFFFF803FFE0FE47FC000070000007C060001F2000C7FE0;
defparam sp_inst_8.INIT_RAM_3A = 256'h0E000001E0000001C0E1C7FFE61FFFFFFFE007FFFFE0038000007000000F8000;
defparam sp_inst_8.INIT_RAM_3B = 256'hFFFE000180080080000004000001E070E1FF9CC3FFFFFFFC0FFFFFF000000000;
defparam sp_inst_8.INIT_RAM_3C = 256'h7FFFFFFFF81FFFFFC00060000000000001800000F078707F81E3FFFFFFFF80FF;
defparam sp_inst_8.INIT_RAM_3D = 256'h7C0C3DFFE0700FFFFFFFFF83FFFFF00004000000000000000000F870787FF00C;
defparam sp_inst_8.INIT_RAM_3E = 256'h0000000170001F073FFFE10E001FFFFFFFE03FFFFF000F000000000000018000;
defparam sp_inst_8.INIT_RAM_3F = 256'hFFFFF807800000000001FC000381FFFFF203F9DBBFFFFFF800FFFFFC01E00000;

SP sp_inst_9 (
    .DO({sp_inst_9_dout_w[30:0],sp_inst_9_dout[10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[10]})
);

defparam sp_inst_9.READ_MODE = 1'b0;
defparam sp_inst_9.WRITE_MODE = 2'b00;
defparam sp_inst_9.BIT_WIDTH = 1;
defparam sp_inst_9.BLK_SEL = 3'b000;
defparam sp_inst_9.RESET_MODE = "SYNC";
defparam sp_inst_9.INIT_RAM_00 = 256'h03FFF80000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0387C000FFDF00000000;
defparam sp_inst_9.INIT_RAM_01 = 256'hFFFFF87FFFC0006FDF80000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC071FC00;
defparam sp_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC0000F0F80000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000F0FC000000FFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_04 = 256'h0007B9C000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000070FC000001;
defparam sp_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFE000007F0C000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sp_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC000007E0600000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000603FFF00001FFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_08 = 256'h00001F0F800079FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000003F9F80003;
defparam sp_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFF8000060603F000E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sp_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80001C0E87F0007FFBFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000F87F001FF83FFFFFFFFF;
defparam sp_inst_9.INIT_RAM_0C = 256'h0060001E0380FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000C0000F81807;
defparam sp_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFC0006000180001E3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sp_inst_9.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFC00030003E02038FF9FFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_0F = 256'h3FE00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0003000CC00061FE0FFFFFFFFF;
defparam sp_inst_9.INIT_RAM_10 = 256'h0000C0E00000021E00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80000003800080;
defparam sp_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFE0000000001804083E01FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0;
defparam sp_inst_9.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80000038001E00203FFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_13 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000078000E00007FFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_14 = 256'h0000008001E001FEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000008001E00;
defparam sp_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFF80000000603C7803FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sp_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFF0FFFFFFFFFFF00000000607C3007FFFFFFFFFFFFFFFFFFFFFFFC;
defparam sp_inst_9.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFE603FFF07FFFFFE000000187810207FFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_18 = 256'h000000018007FFFFFFFFFFFFFFFFFFFFFFF8007FC01FFFFFFC0000001018003F;
defparam sp_inst_9.INIT_RAM_19 = 256'hF000FFFFFFF8000000080E00FFFFFFFFFFFFFFFFFFFFFFFF000FE003FFFFFF80;
defparam sp_inst_9.INIT_RAM_1A = 256'hFFFFFFFFF80070003FFFFFFE0000000000E01FFFFFFFFFFFFFFFFFFFFFFFE003;
defparam sp_inst_9.INIT_RAM_1B = 256'hFFFFFFFFFFFFF8FFFFFFFE000C0007FFFFFFC0000000000403FFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_1C = 256'h00000000018FFFFFFFFFFFFFFF0FFFFFFFC0400001FFFFFFF80000000020007F;
defparam sp_inst_9.INIT_RAM_1D = 256'h000FFFFFFFE000000000000FFFFFFFFFFFFFFFF0FFFFFFF81C00003FFFFFFF00;
defparam sp_inst_9.INIT_RAM_1E = 256'hF87FFFFFC3F80003FFFFFFFC000000000000FFFFFFFFFFFFFFFF87FFFFFE0FC0;
defparam sp_inst_9.INIT_RAM_1F = 256'hFFFFFFFC07FFFFC3FFFFF87F0000FFFFFFFF8000000000000FFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_20 = 256'h00000000001FFFFFFFFF0001FFF81FFFFF0FE0007FFFFFFFE0000000000060FF;
defparam sp_inst_9.INIT_RAM_21 = 256'h07FFFFFFFF80000000000003FFFFFFFFF00000FF83FFFFE1FC001FFFFFFFFC00;
defparam sp_inst_9.INIT_RAM_22 = 256'hFF07FFFFCFF003FFFFFFFFF00000000000007FFFFFFFFF00000FF87FFFFE7F80;
defparam sp_inst_9.INIT_RAM_23 = 256'hFFFFFFFFC0000FF0FFFFF1FC01FFFFFFFFFE0000000000000FFFFFFFFFF80000;
defparam sp_inst_9.INIT_RAM_24 = 256'h00000000003FFFFFFFFFFE0001FF1FFFFE3F83FFFFFFFFFFE0000000000001FF;
defparam sp_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFF00000000000007FFFFFFFFFFE0001FE3FFFFE7F3FFFFFFFFFFF800;
defparam sp_inst_9.INIT_RAM_26 = 256'hBFC7F3FF9FBFFFFFFFFFFFFC000000000000FFFFFFFFFFFF8001FC7FFFFCFFFF;
defparam sp_inst_9.INIT_RAM_27 = 256'hFFFFFFFFFFF9FFF9FFFFFFF7FFFFFFFFFFFFC000000000001FFFFFFFFFFFFC01;
defparam sp_inst_9.INIT_RAM_28 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC000000000003FF;
defparam sp_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFF9800E00000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC0;
defparam sp_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFE393C000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC7F10000000003FFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_2C = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFE00000000007FF;
defparam sp_inst_9.INIT_RAM_2D = 256'hFFFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sp_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFE000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFFFF8000000000007FFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_30 = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFC7FFFFFFFFFFFFE000000000000FFF;
defparam sp_inst_9.INIT_RAM_31 = 256'hFFFFFFFFFF0000000000003FFFFFFFFFFFFFFFFFFFFFFFF8FFFFFFFFFFFFFC00;
defparam sp_inst_9.INIT_RAM_32 = 256'hFFFFFFFFF0FFFFFFFFFFFFE0000000000007FFFFFFFFFFFFFFFFFFFFFFFF8FFF;
defparam sp_inst_9.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFC1FFFFFFFFFFFF8000000000000FFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_34 = 256'h0000000003FFFFFFFFFFFFFFFFCFFFFFFF87FFFFFFFFFFE00000000000001FFF;
defparam sp_inst_9.INIT_RAM_35 = 256'hFFFFFFFF800000000000007FFFFFFFFFFFFFFFF9FFFFFFF0FFFFFFFFFFF80000;
defparam sp_inst_9.INIT_RAM_36 = 256'hE3FFFFFF87FFFFFFF9FFF00000000000000FFFFFFFFFFFFFFFFF1FFFFFFE1FFF;
defparam sp_inst_9.INIT_RAM_37 = 256'hFFFFFFFFFFFFFC3FFFFFF0FFFFFFFC7FFC00000000000001FFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_38 = 256'h0000000007FFFFFFFFFFFFFFFFC7FFFFFE1FFFFFFC3FFF800000000000003FFF;
defparam sp_inst_9.INIT_RAM_39 = 256'hFF9FFCF8000000000000007FFFFFFFFFFFFFFFF8FFFFFF83FFFFFE0FFFF00000;
defparam sp_inst_9.INIT_RAM_3A = 256'hF1FFFFFE1FFFFFFFFF1E000000000000001FFFFFFFFFFFFFFFFF8FFFFFF07FFF;
defparam sp_inst_9.INIT_RAM_3B = 256'hFFFFFFFFFFFFFF7FFFFFFBFFFFFFFF8F0000000000000003FFFFFFFFFFFFFFFF;
defparam sp_inst_9.INIT_RAM_3C = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFE7FFFFFFF8780000000000000007FFF;
defparam sp_inst_9.INIT_RAM_3D = 256'hFFF3C000000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F80000000;
defparam sp_inst_9.INIT_RAM_3E = 256'hFFFFFFFE8FFFFFF8C000000000000000001FFFFFFFFFFFFFFFFFFFFFFFFE7FFF;
defparam sp_inst_9.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFE03FFFFFE00000000000000000007FFFFFFFFFFFFFFFF;

SP sp_inst_10 (
    .DO({sp_inst_10_dout_w[30:0],sp_inst_10_dout[11]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11]})
);

defparam sp_inst_10.READ_MODE = 1'b0;
defparam sp_inst_10.WRITE_MODE = 2'b00;
defparam sp_inst_10.BIT_WIDTH = 1;
defparam sp_inst_10.BLK_SEL = 3'b000;
defparam sp_inst_10.RESET_MODE = "SYNC";
defparam sp_inst_10.INIT_RAM_00 = 256'h6230F95C3FFFF82C20182FF4CDFFB41130F18E3FF7FE8B3E5AEA4F0763E1FFFF;
defparam sp_inst_10.INIT_RAM_01 = 256'h77EFC6B827DF4B0107FDC7FFFCFE781C847FD93FC0021E3E31C3FE3F76B9DE3E;
defparam sp_inst_10.INIT_RAM_02 = 256'h7E003D8C00840FE5FC4E920974AEA03C28FFFFEF81D9DE83F803F0006BCFCC30;
defparam sp_inst_10.INIT_RAM_03 = 256'h07FC46CC67E403C01FC0D01181FD8FA2F3E74BADAE40DE8FFFF0000C67EF7E20;
defparam sp_inst_10.INIT_RAM_04 = 256'hEE4700173FFFFE8475A80E7C00BC0FFC0823F07F20AC9FCF9367896005F0FFFE;
defparam sp_inst_10.INIT_RAM_05 = 256'hF9E9140184CF6DEED8210FFFFFC1FB3EB8672013C7DFE184C423CFC7D8386A0C;
defparam sp_inst_10.INIT_RAM_06 = 256'h9FF9FFE39218FF39E5800A423C347F840E7FFFC3F1F22B84000E7FCBFE1CF007;
defparam sp_inst_10.INIT_RAM_07 = 256'hA9401007FC0013807FFEE0431E467F9E00F5315E6DB80375FFF09C07E37EC001;
defparam sp_inst_10.INIT_RAM_08 = 256'h68EF806010FFA148D65CFF6031F09E0C1E08FFC89FE3F80E91D3DD3D90222FFD;
defparam sp_inst_10.INIT_RAM_09 = 256'h38FFC21A1B4DCA3A6B0F82F7FB4082BC0FE0066E3D99BBF11FF1C7FE3380D050;
defparam sp_inst_10.INIT_RAM_0A = 256'hD98931270BA00303F803E77673F4F61030F8BF019573E1FC18CCCF87B93C17C6;
defparam sp_inst_10.INIT_RAM_0B = 256'hB2C187C22181B9BDE610626003F87FC01FE930CACB5870025BEBDB947E3B811D;
defparam sp_inst_10.INIT_RAM_0C = 256'h12FC472DFC51C093ED38403873B23C520C59C0770FFC01FD15834320980384D8;
defparam sp_inst_10.INIT_RAM_0D = 256'h24607FE0F3889191F8F97D3E25EB873328079F7C4402239B783863E3F03FBF78;
defparam sp_inst_10.INIT_RAM_0E = 256'h2E5C0C1E17F3A288DFFF0C1073FD0FF07DEDEB2C70B82C867963182134F20F1F;
defparam sp_inst_10.INIT_RAM_0F = 256'hA65805B3EE70019F01C371BA74527BFCF982FACCC27D8CA7FF7064E30D987F10;
defparam sp_inst_10.INIT_RAM_10 = 256'h278F4FA2A06CE8813C371EC60039E4F84C262EABE67FBF80549E1EC2A8970336;
defparam sp_inst_10.INIT_RAM_11 = 256'hD1FF66079957C1B6B37A3678AAAC93A5B9CC800CA4DE0A02C3F7BE1E7DF04C2F;
defparam sp_inst_10.INIT_RAM_12 = 256'hA096DE6A3128366CEF3C780659EDE4D10B415B24878279FC93E1849CFB40D96C;
defparam sp_inst_10.INIT_RAM_13 = 256'h9BF6C303BC96FDCAEA8CBC8E0C9C3EF04F00F5C73FD2B458D1958E33E91FDE8F;
defparam sp_inst_10.INIT_RAM_14 = 256'hDE049CCE5D3D729454F1FBB5F3BF6ED1871B7F70973C687F2626803557F6137A;
defparam sp_inst_10.INIT_RAM_15 = 256'h625AF80FDF9C396760D17241BDC84ABE1FC2B008ECF261E9442495AAC60FFCF8;
defparam sp_inst_10.INIT_RAM_16 = 256'h71913E9159904C6DBF5FF3F44236F01ABBDF1C56964F638015A19D9F1CEF376B;
defparam sp_inst_10.INIT_RAM_17 = 256'hDC04183C60DC7802A7E48F111D456650783F6B00C66A74C56C0BAECFE3E002BA;
defparam sp_inst_10.INIT_RAM_18 = 256'h18673796DDFD67FE60099F1CBC4010431DD33F5E4CA0CC03FAC3C4BB8971AB68;
defparam sp_inst_10.INIT_RAM_19 = 256'hAB0BFE500F1D46EA7E9504FC27FE3800C361BE3F871747A5D872F318BB00785C;
defparam sp_inst_10.INIT_RAM_1A = 256'h3E8DE17D750E1B6E924E07F8A1CFE47CCC4813F79E000CFF39B809E72BF9543B;
defparam sp_inst_10.INIT_RAM_1B = 256'h0CE18E12384228F1DC0E4B4629B82AFA60FA47B86F32B2C94E387787FF0AC7D2;
defparam sp_inst_10.INIT_RAM_1C = 256'h7898A704C7560138661B500B8D258649C1276E8181DA0F9FE81787CE744EC45C;
defparam sp_inst_10.INIT_RAM_1D = 256'hB4E6C13E3F9728C139FC3498C0DF3CC6FDFB7B563ECEE09312022A66E0F3F5D3;
defparam sp_inst_10.INIT_RAM_1E = 256'hA8741C392139D650A2C7C7D6FFD87FC681EF9C3BE78FDE0B05E30259D97B32D8;
defparam sp_inst_10.INIT_RAM_1F = 256'h1F8FF0E9E71B3A8170862413F689007878E0EFF11A7E72B573877C7F0A10E321;
defparam sp_inst_10.INIT_RAM_20 = 256'hCE46C0F09ED807C1FF968B4DEBAB95CF9C82780440BF070135A5633F346E6BE0;
defparam sp_inst_10.INIT_RAM_21 = 256'h5704007E0A1D0D891929BFFDE3E01E4B8B49AE3AAB2267178970A0A003F01713;
defparam sp_inst_10.INIT_RAM_22 = 256'hBB76BE21499B7C6900078FDA010DE53819DFB1F803FCB842CCCBA4B4F4EE7D42;
defparam sp_inst_10.INIT_RAM_23 = 256'h00C3E1DB681BC3969F3DEC2F2E68A00837B8CE19FF9CB86575FE207F2B9A5CB3;
defparam sp_inst_10.INIT_RAM_24 = 256'h0980639C7237F1047FE2C513747DD06725C5CEB4A1008CFFD39B98F7EE7EEDBF;
defparam sp_inst_10.INIT_RAM_25 = 256'h478EFFC67EEC030702236F637F400FF9444400576B2C40F8188A287F3F9FE720;
defparam sp_inst_10.INIT_RAM_26 = 256'h6600119E6670FAD415F3B8231B162F6DE8F323E0038C6B1AFA2E7024763B2DF6;
defparam sp_inst_10.INIT_RAM_27 = 256'hCC19E9DED94924D97C2CE8C8DE4C447C391B9696F167FE9E567C20649D533522;
defparam sp_inst_10.INIT_RAM_28 = 256'hCEDB0E71FFD3FF093C1E5B0C02C2BA1B0449259B890F80331FE036357BC6FECF;
defparam sp_inst_10.INIT_RAM_29 = 256'h0C0EF80E7749A0DBA35446E27FE3A7F817D3FD361F87488C0C0F6A43E067E01B;
defparam sp_inst_10.INIT_RAM_2A = 256'h821C97532D35C1A1E00784BEC9AC1C6180FBC7FE242207B247FCF17F3610C24E;
defparam sp_inst_10.INIT_RAM_2B = 256'hF19CC0F8F8219A0F14189038B8062C031C20570E5983808EF07FBC8C39E40CEC;
defparam sp_inst_10.INIT_RAM_2C = 256'h80665DB9FA9FFC30E006279A240199BFFEC5AFE2899F18757BDB67F86BD02807;
defparam sp_inst_10.INIT_RAM_2D = 256'hEF2005BF891F820C01BEF353FF0E0E3FFCFB9C63E2FCED40D5F3D639A1474D6D;
defparam sp_inst_10.INIT_RAM_2E = 256'h75D9EDCCF8658FBC408C20F5CE27E1019FBA7F03F00EC01F61E54E23CD870ABC;
defparam sp_inst_10.INIT_RAM_2F = 256'h0EE07FE0213434FDC041BB801E6FB0FFFBB8D39F8FFB7D1647E07E03C800313A;
defparam sp_inst_10.INIT_RAM_30 = 256'h40071F196CCFC1FF0FC040CCF43EBF005CC88F12172FE2BB6642003FB7EBE87C;
defparam sp_inst_10.INIT_RAM_31 = 256'hE7BF884AB50B9C00E36A1388FC1FF000063F9FC7B26E6CD4F08F19CCD8152E54;
defparam sp_inst_10.INIT_RAM_32 = 256'h2CE3C002DF427FE20173C7980D800EFA38710FF7FF0E03E1C7B3354EC42EA233;
defparam sp_inst_10.INIT_RAM_33 = 256'hC27E40F003DDF61CF0B079E701F41003E95E41C001809FFF70FE7FF1F800279D;
defparam sp_inst_10.INIT_RAM_34 = 256'h00CA06DFF331FC03901E306F82F3983F8710E0617D0EF0341F99041606EF878F;
defparam sp_inst_10.INIT_RAM_35 = 256'hFC7D8DC220C3300425C47F123FE0000FC40AC1E6B327F0D329894833AE7BBD33;
defparam sp_inst_10.INIT_RAM_36 = 256'h1CEEC004B2BF74BF2666D1838B90797D81D56F7E7FCF180180F8E67E7E2BA4B1;
defparam sp_inst_10.INIT_RAM_37 = 256'hFB3FFF001FFE6C7BAC10BE13978869528CC1FBF01F4B19A0B67FD9F3FF81FFF9;
defparam sp_inst_10.INIT_RAM_38 = 256'h90C70E4781260F9CFFC00061DC08CFC0974B79BE56ED26A87F60827E11A65A67;
defparam sp_inst_10.INIT_RAM_39 = 256'hC7D6B36DB130082915F1E2E64039F83FE038B8CD20F000A770D8F65C05CE1F81;
defparam sp_inst_10.INIT_RAM_3A = 256'h8AC3B0C4A34D7B0FD6D6D32400C8298B8856F9C0003FFE7FFF8EF45E96342BD3;
defparam sp_inst_10.INIT_RAM_3B = 256'h7FE3001FE0FC6EAC0618B8633F491E467E4D001852607FE26BFE0C087CFE67F1;
defparam sp_inst_10.INIT_RAM_3C = 256'hF031348698A4601E6620FBA20624861816141992F20C8432BC0C33EA732B2340;
defparam sp_inst_10.INIT_RAM_3D = 256'h0A0C3DE0C4073477060D6214F87FCE931FE70078917D82770FE5F398B81A6431;
defparam sp_inst_10.INIT_RAM_3E = 256'hFF21E4279E0C968CF53FCC60308CFC49EF5687E7F1A49F3CF31FDB2F906F51D1;
defparam sp_inst_10.INIT_RAM_3F = 256'h10F1E8AF3FBB87ECB7997DE16BD858A2E0DC67805F3CB366CC06380579E61C3F;

SP sp_inst_11 (
    .DO({sp_inst_11_dout_w[30:0],sp_inst_11_dout[12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[12]})
);

defparam sp_inst_11.READ_MODE = 1'b0;
defparam sp_inst_11.WRITE_MODE = 2'b00;
defparam sp_inst_11.BIT_WIDTH = 1;
defparam sp_inst_11.BLK_SEL = 3'b000;
defparam sp_inst_11.RESET_MODE = "SYNC";
defparam sp_inst_11.INIT_RAM_00 = 256'h1E3FFD6000001FD01FF8100BF3FFB41F30F18FC007FDF9C2B319CFFFB4000000;
defparam sp_inst_11.INIT_RAM_01 = 256'h880FEA7C46C8B2F1FFD6000003FF87E383803EFFC003FE3E31FC003FDE486942;
defparam sp_inst_11.INIT_RAM_02 = 256'hFE003E7C0087F019F9A708279EE1BFFEB000001FFE063E7C07FFF00077CFCC3F;
defparam sp_inst_11.INIT_RAM_03 = 256'hFFFF81CC181BFBC01FFFC011FE020F260004EE339FBFEB00000FFFF01FE081DF;
defparam sp_inst_11.INIT_RAM_04 = 256'h1FDFFFE20000018079980183FFBC0FFFF823FF80C0B27FF0827878FFFEA00001;
defparam sp_inst_11.INIT_RAM_05 = 256'h06100C01F9AFB3E05FDE500007DFFBBD8018DFF3C7DFFF84FFDC3007B83F8017;
defparam sp_inst_11.INIT_RAM_06 = 256'h9FFFFFFF93E700C603800F91F9F3B7FBF48000C7FFFC1803FFFE7FFBFFFCFFF8;
defparam sp_inst_11.INIT_RAM_07 = 256'hC73FF00003FFF3FFFFFFE07CE039807E00F8E39EF77FFFA6001063FFFF003FFF;
defparam sp_inst_11.INIT_RAM_08 = 256'hF0F87F9FE5004A3F0FC0009FCFFF7FFFFE0F0007601FF80F34CCC1FBFFFCB003;
defparam sp_inst_11.INIT_RAM_09 = 256'h07003FFA1D9D27BEF0F07F580C9F01BC001FF9EFC3E7C7F1E0003801FF80E53E;
defparam sp_inst_11.INIT_RAM_0A = 256'hDE060E1F0C0000FC07FFE7BA3CB8D4CFCFF2C1561B13E003FF3CF07870FC2800;
defparam sp_inst_11.INIT_RAM_0B = 256'h21C19FC1DFFE79C001CFE3800387803FFFF188F9E865FFFF8C081C73FE047FE3;
defparam sp_inst_11.INIT_RAM_0C = 256'h1FF7C71E039A17B00CF83FFF8FBC0039FC61C070F003FFFE1303D23F87FC7965;
defparam sp_inst_11.INIT_RAM_0D = 256'hE380001FFC2511F978FB82C0B3A7800F07FFE0FF80077F9C783E1C000FFFC2D0;
defparam sp_inst_11.INIT_RAM_0E = 256'hF05C13FE7BF3BE70C000FFE523FF4BFF3E120ECBFF87E07FFE9FE020CFF3CF1F;
defparam sp_inst_11.INIT_RAM_0F = 256'h66E013801E7FFE5F027F7F3E77CC780307FCA8FCF6BE5FC0005A1F1F7C07FFEF;
defparam sp_inst_11.INIT_RAM_10 = 256'h078E6EB6401385323D7001C7FFC1E00FCFF7EED80600407F9A5E1FBCDC8800C6;
defparam sp_inst_11.INIT_RAM_11 = 256'h360098007E90C1F0EF83F18063FA200C403CFFF03C01FBFCFFF98001800FF09B;
defparam sp_inst_11.INIT_RAM_12 = 256'h40F547EDC1DFC293103C07FA59FC0445F73E4077E78106039C1E07803F7F1EFF;
defparam sp_inst_11.INIT_RAM_13 = 256'hD971C0FC03E601CE89FCC031F043C0FFC0FF79FF0010DFC1E089F20FE6E03F00;
defparam sp_inst_11.INIT_RAM_14 = 256'h3E031DEE232349B7CC0E0079F03FE03F880C006878201800CEB9800935F15218;
defparam sp_inst_11.INIT_RAM_15 = 256'hA19CF400003DC6E700C9767FF4987981E03F3E0FFC0FE009803D8E33DE0001EF;
defparam sp_inst_11.INIT_RAM_16 = 256'h7FF007987DFF540E3D200004FDCEF002D3454E3A66C09C7FE661FF80FCC3276C;
defparam sp_inst_11.INIT_RAM_17 = 256'h3C03E7C3FF10FFFE80E70FAE1EC67A8F80003FFFC669BC83BA069F201C1FFCC6;
defparam sp_inst_11.INIT_RAM_18 = 256'hC7FFF01EEE04E001FFFE7FE10FBFD03FE1E43F7F6EBBF0001C1C3CFFB3258CE6;
defparam sp_inst_11.INIT_RAM_19 = 256'h3255AF900075B91DFE09D083E001FFFFFF7E21C07F10F8391FE725B97C0003E7;
defparam sp_inst_11.INIT_RAM_1A = 256'h3E7CE38199FE53D0A66E00083E301C7C0E0FF0087FFFFFFFC24007E71C0E67F8;
defparam sp_inst_11.INIT_RAM_1B = 256'hF3FE0011FF85CFEFDC70727E252B13F3E00467C780F3816A7E078FF800FEF86C;
defparam sp_inst_11.INIT_RAM_1C = 256'h876067001A61FEFF861CCFF3F9DC7FC6064F0ED4F3BCFF802C18780270363843;
defparam sp_inst_11.INIT_RAM_1D = 256'hE725EEFE009737FE07FC08B43F3FC0C704047F99E1FE00DB0DE82F0F7FF00593;
defparam sp_inst_11.INIT_RAM_1E = 256'hCFF3FC3E430D2C897B3FC00EFFFF803F800F43C7F80061FB07FDFE3FC1722EA1;
defparam sp_inst_11.INIT_RAM_1F = 256'hFFF00F321F00FCFF0F87C84D49995E87F8044FFFE181F0826078FF80F3E01FDF;
defparam sp_inst_11.INIT_RAM_20 = 256'hFF8031F10107FFFE007A4743E7CC70FFE109A7FC9720FF0189A6FC000C00F31F;
defparam sp_inst_11.INIT_RAM_21 = 256'h6577FFFE021DFFF0E61F80001FFFE187C938617CC71DF825757F75CFFFF01007;
defparam sp_inst_11.INIT_RAM_22 = 256'hFD8E41C183CBD6DDFFFF805BFFF21EC7F8200FFFFC007C31C42FC8730F0C2EE3;
defparam sp_inst_11.INIT_RAM_23 = 256'hFFFC1E3D5DF867D98001F17425273FF7F0480FFE0063C7E203FFDF80C7C9226F;
defparam sp_inst_11.INIT_RAM_24 = 256'hEE7F8062700FFEFF8001EEFF05F93000262EA1933FFFFC013DE7E708118E027F;
defparam sp_inst_11.INIT_RAM_25 = 256'hFB8EFFC1864FFFFFFC1CCF00FFBFF001DE91403FB72000C5D279CFFFFF80223F;
defparam sp_inst_11.INIT_RAM_26 = 256'hBF781F9F9095FCD01DF0476A1FF6314219F71FFFFC0076ECAC18FBE4763C9651;
defparam sp_inst_11.INIT_RAM_27 = 256'hFFE1E1E1C18F0DEF7FE0F6147F8007FC00E9C0F0FF0801FE31FFFF841E302639;
defparam sp_inst_11.INIT_RAM_28 = 256'h005E000FFFCFFFFE3C1F870FFCDCFE1807C2ABE001FF800D5A003DC6003FFA3F;
defparam sp_inst_11.INIT_RAM_29 = 256'h000FF80E0498C213C00FC0E1FFFFC7F8183001DD9FB800FC7D70087FE0602BF4;
defparam sp_inst_11.INIT_RAM_2A = 256'h001C78E3DE8C0021E007808E2831F00FF0183FFFF823FFBE3FB9C170C11FCE20;
defparam sp_inst_11.INIT_RAM_2B = 256'hFFE0C0F8001EE40F0FFF1FD780063C03FC315E0B8601FE020FFFFF0C3FE403F7;
defparam sp_inst_11.INIT_RAM_2C = 256'h7F804679FB7FFFFF00061819CA4187FFF3FC60038F9FE7F7144FF80031C017FF;
defparam sp_inst_11.INIT_RAM_2D = 256'hE1FFF980729E7FF0007EFF6FFFFFF1C0030381CBE1FCEE7FCC03C7FFC0FFA826;
defparam sp_inst_11.INIT_RAM_2E = 256'h67C9FDF487220C3FBF001E95BFF800099FBDFFFFFFF03FE060317E63CDC4F980;
defparam sp_inst_11.INIT_RAM_2F = 256'hFEFF801FFE303EFBFFFEBC68E00FCF00079C6FE000017DC7BFFFFFFC07FFC102;
defparam sp_inst_11.INIT_RAM_30 = 256'h80000FFF0C3FFFFFF03FBF0007DE7FFF9C85801218C006D40A7C00007FF867FF;
defparam sp_inst_11.INIT_RAM_31 = 256'hE7C007F3163C60000177F387FFFFFFFFFFC0007B8FF1F0D8500F1A3027E56DDB;
defparam sp_inst_11.INIT_RAM_32 = 256'hCE1FFFFCEE407FF000E08E23F000003BBFF0FFFFFFFFFFFE004432FF3FCF2A03;
defparam sp_inst_11.INIT_RAM_33 = 256'hFFFFFF0FFC1C7BC3FF7FBDCF01F81F6008A63E00007FFFFF0FFFFFFFFFFFC001;
defparam sp_inst_11.INIT_RAM_34 = 256'h0009FFFFF30FFFFFFFE1CF8F83487FFFF7B5E07E7E8E009CA061000FFFEF807F;
defparam sp_inst_11.INIT_RAM_35 = 256'h01907366AB0000001BFC7FF1FFFFFFF03BF3C0498FFFFEE6998E8FF26053AE0C;
defparam sp_inst_11.INIT_RAM_36 = 256'hA21FBFF9367F48C936B7A0000810063D8F031F7F803007FE000D11FFFFCD93B1;
defparam sp_inst_11.INIT_RAM_37 = 256'hFC0000FFE0007627D3EF2E8FF808328CD0A00380008719E071FFE00C007E0001;
defparam sp_inst_11.INIT_RAM_38 = 256'h8038F104F8E1FFE0003FFF801F45F03FE5D8FE001AB6312000600181F1A7861F;
defparam sp_inst_11.INIT_RAM_39 = 256'h1E9938EB00C0081E0E10385E3FFE07C01FC080E89F07FEBD10972D5B0FFC0001;
defparam sp_inst_11.INIT_RAM_3A = 256'hE03C0F38A8F1C3C59B54147800C7C7F78F1207FFFFC00180000CA3E069D767E6;
defparam sp_inst_11.INIT_RAM_3B = 256'h7FFC000000007D63E1E7011C301528EF1EFE00198DFFFFE227FFFFF000000001;
defparam sp_inst_11.INIT_RAM_3C = 256'h800EFFFE059C601F87E0002007FC7867E43BE011F52494133C0C0005FFE366C0;
defparam sp_inst_11.INIT_RAM_3D = 256'h8C9258E084073000FFF2E0B3F87FF7700007007D8E827C82F003FB48AB438431;
defparam sp_inst_11.INIT_RAM_3E = 256'hF71E1BC43FF1B71ECBE08C60308003D61F327FE7FE3B8000F31FB8D06FB17E20;
defparam sp_inst_11.INIT_RAM_3F = 256'hF0FE129BBFC786E3C86278FE6783FF7B00DC060040CBFD6643FE3FF984001FFF;

SP sp_inst_12 (
    .DO({sp_inst_12_dout_w[30:0],sp_inst_12_dout[13]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13]})
);

defparam sp_inst_12.READ_MODE = 1'b0;
defparam sp_inst_12.WRITE_MODE = 2'b00;
defparam sp_inst_12.BIT_WIDTH = 1;
defparam sp_inst_12.BLK_SEL = 3'b000;
defparam sp_inst_12.RESET_MODE = "SYNC";
defparam sp_inst_12.INIT_RAM_00 = 256'h01C0018000001FFFFFF8000000004BE0CF0E700007FEF84923F8300038000000;
defparam sp_inst_12.INIT_RAM_01 = 256'h000FF200276F820E0018000003FFFFFF800000003FFC01C1CE00003F9E0EF27E;
defparam sp_inst_12.INIT_RAM_02 = 256'h01FFC003FF780001FE1FF835F0E04000C000007FFFFFFE0000000FFF803033C0;
defparam sp_inst_12.INIT_RAM_03 = 256'hFFFFFFCC0000043FE0003FEE00000FDE00068E3F80000C00000FFFFFFFE00000;
defparam sp_inst_12.INIT_RAM_04 = 256'hFFC0000400003F807E7800000043F00007DC000000BE0000DC7FF80000C00001;
defparam sp_inst_12.INIT_RAM_05 = 256'h000003FE01303FE020006000003FFBC38000000C3820007B0000000787C00BE7;
defparam sp_inst_12.INIT_RAM_06 = 256'h600000006C000000007FF01A01F030000700003FFFFFF8000001800400030000;
defparam sp_inst_12.INIT_RAM_07 = 256'h00FFF00000000C0000001F8000000001FF01401E07000038000FFFFFFF000000;
defparam sp_inst_12.INIT_RAM_08 = 256'h00F8000006000EFFFFC000000000000001F00000000007F026C0C1F80000C000;
defparam sp_inst_12.INIT_RAM_09 = 256'h00000005E1E9E03E000000600FBFFFBC000000100000000E00000000007F065E;
defparam sp_inst_12.INIT_RAM_0A = 256'h20000000F00000000000183CBF80C8C0000300CFE0F3E000000300000003C000;
defparam sp_inst_12.INIT_RAM_0B = 256'hC03E7FC00000060000001C00038000000001D0F8087C00001027E00FFE000000;
defparam sp_inst_12.INIT_RAM_0C = 256'h1E07C700001CE78FF3F80000004000000381C070000000001A03CC3F80000183;
defparam sp_inst_12.INIT_RAM_0D = 256'hE0000000003611F678F80000DA607FFF0000000000000060783E000000000360;
defparam sp_inst_12.INIT_RAM_0E = 256'h005C000183F3BE00C000000643FF33FF00000C98007FE00000000020000C0F1F;
defparam sp_inst_12.INIT_RAM_0F = 256'hE6000F800180001F0000803E77C078000000CCFCF13FC00000660000FC000000;
defparam sp_inst_12.INIT_RAM_10 = 256'h078E8E4600007DEC3CF000380001E0003007EEF8060000001C9E1F80FB000009;
defparam sp_inst_12.INIT_RAM_11 = 256'hF0000000001AC1F0E003F0001DC5C01C000300003C000400FFFF8000000000D3;
defparam sp_inst_12.INIT_RAM_12 = 256'h00F4401001FFFE00003C000319FC0439FF0047F8587F00006000078000801FFF;
defparam sp_inst_12.INIT_RAM_13 = 256'h270FC000000601CE8803003FFFC000FFC00051FF00171FC0007E09FFE0000000;
defparam sp_inst_12.INIT_RAM_14 = 256'hFE001C0E00C087883C000001F03FE000700FFF98003FF8000B3F800109F04C07;
defparam sp_inst_12.INIT_RAM_15 = 256'h601F0C000029FFE700C671800447878000003E0FFC001E09FFC3803C3E00014F;
defparam sp_inst_12.INIT_RAM_16 = 256'h7FF000607E004C0FC30000067FFEF00263393009F9C0000007E1FF8003033890;
defparam sp_inst_12.INIT_RAM_17 = 256'hFC000000001FFFFE80180FC01DC7824000006FFFC668330039FE7FE0000000FE;
defparam sp_inst_12.INIT_RAM_18 = 256'hFFFFF01D0FFBE00000000001FFFFD00001F83F3F8F680000141FFCFF83198FE1;
defparam sp_inst_12.INIT_RAM_19 = 256'hC39D60100059FFFFFE01CEFFE000000000803FFFFF10003E1FEFC63300000287;
defparam sp_inst_12.INIT_RAM_1A = 256'hC1FCE001E1FE239FD18E000D3FFFFC7C0EEFF0000000000003FFFFE7000F87F9;
defparam sp_inst_12.INIT_RAM_1B = 256'h000000100007F01FDC007C7E21CCE603E000C7FFFFF380647E0000000001007F;
defparam sp_inst_12.INIT_RAM_1C = 256'hFFFFE70019800000061FC003FE03FFC0078F0EE60A80FF80381FFFFE70060040;
defparam sp_inst_12.INIT_RAM_1D = 256'h184C0FFE00C73FFFFFFC008E000000C7FC007FE01FFE00E301F3D1A07FF00713;
defparam sp_inst_12.INIT_RAM_1E = 256'hF00FFC3F80F6431303FFC014FFFFFFFF800EC00000007FFB07FE01FFC17C213D;
defparam sp_inst_12.INIT_RAM_1F = 256'h0000003C00FFFF00FF87F03E9063C0FFF8068FFFFFFFF0806800000003FFFFFF;
defparam sp_inst_12.INIT_RAM_20 = 256'hFFFFFFF00000000000037F401FF00FFFFE07D402B03FFF01D1A7FFFFFC000300;
defparam sp_inst_12.INIT_RAM_21 = 256'hD307FFFE035DFFFFFFFF8000000000001D07E0FF00FFFFC4FB80AC0FFFF01A07;
defparam sp_inst_12.INIT_RAM_22 = 256'h7E01FFFE07E3CDC1FFFF8073FFFFFFFFF80000000000015FC3E7F00FFFF01F3C;
defparam sp_inst_12.INIT_RAM_23 = 256'h000000019607CFE07FFE00F9DCE03FFFF00D0FFFFFFFFFE000000000001241E1;
defparam sp_inst_12.INIT_RAM_24 = 256'hEFFFFFFE70000000000008A0FEFE0FFFD81F20703FFFFC01A1FFFFFFFFFE0000;
defparam sp_inst_12.INIT_RAM_25 = 256'h038EFFC0048FFFFFFFFFCF0000000001C0E67FAFC0DFFF03E1F80FFFFF80343F;
defparam sp_inst_12.INIT_RAM_26 = 256'h1F87E0600F0C00D01DF0004C1FF63F7FF9F0000000007E0F3005FC1B89C07830;
defparam sp_inst_12.INIT_RAM_27 = 256'h0001E1FFC1F0F3F0801F01E3C00007FC000DE0F0FF0FFFFE100000041FF03838;
defparam sp_inst_12.INIT_RAM_28 = 256'h0023FFFFFFC000003C1FFF0FFF3F01E7F83C580001FF80019C003C07FFFFFA00;
defparam sp_inst_12.INIT_RAM_29 = 256'h000FF80E06FC01E3FFFFC0E0000007F81FF001E3E07FFF038300087FE06033D0;
defparam sp_inst_12.INIT_RAM_2A = 256'hFFE3FFFC007C0021E00780D297C1FFFFF01800000023FFBE003E3E8FFFE031E0;
defparam sp_inst_12.INIT_RAM_2B = 256'h0000C0F80000FFF0FFFFE00F80063C03FC3ADFF3FFFFFE020000000C3FE40007;
defparam sp_inst_12.INIT_RAM_2C = 256'hFFFFBFF9FB000000000600180E7E7FFFFC03E0038F9FFFF6706FFFFFFFC00000;
defparam sp_inst_12.INIT_RAM_2D = 256'hE1FFFE7FFC6BFFFFFFFEFF6000000000000381CC1FFCEF803C03C7FFFFFFCBB7;
defparam sp_inst_12.INIT_RAM_2E = 256'h7839FDFB00E00C3FFFFFFF08FFFFFFF99FBC000000000000603181E3CDF80780;
defparam sp_inst_12.INIT_RAM_2F = 256'h0100000000303F07FFFF4018000FFFFFFFDB3FFFFFFF7DC78000000000000102;
defparam sp_inst_12.INIT_RAM_30 = 256'hFFFFFFFF0C0000000000000007E1FFFFE30380121FFFFEE6DE7FFFFFFFF86000;
defparam sp_inst_12.INIT_RAM_31 = 256'hE7FFFFFC08BFFFFFFF7FF380000000000000007C7FFFFF20300F1BFFFFF915DF;
defparam sp_inst_12.INIT_RAM_32 = 256'hF1FFFFFF0EC07FFFFFFF002FFFFFFFFBBFF00000000000000007CFFFFFF02603;
defparam sp_inst_12.INIT_RAM_33 = 256'h00000000001C7C3FFFFFC1DF01FFE0FFF6FBFFFFFFFFFFFF0000000000000001;
defparam sp_inst_12.INIT_RAM_34 = 256'hFFF7FFFFF30000000000000F8387FFFFF833E07F8071FF233FFEFFFFFFEF8000;
defparam sp_inst_12.INIT_RAM_35 = 256'hFE0E00F6D3FFFFFFFFFC7FF0000000000003C0707FFFFF06798FF00C1F9C4FFF;
defparam sp_inst_12.INIT_RAM_36 = 256'hC1FFFFFE31FF7F06C678FEFFF7EFFFFD8F0F008000000000000E0FFFFFF18FB1;
defparam sp_inst_12.INIT_RAM_37 = 256'h000000000000781FFFFFCE7FFFF7C3BF1F3FFC7FFFFF19E1F000000000000001;
defparam sp_inst_12.INIT_RAM_38 = 256'h7FFFFF04FFE00000000000001F83FFFFF9C7FFFFE36FC7CFFF9FFFFFF1A7FE00;
defparam sp_inst_12.INIT_RAM_39 = 256'hE0F7C3EDFFFFF7FFFFF0383E00000000000080F07FFFFF3CF0EFC1B7F7F7FFFE;
defparam sp_inst_12.INIT_RAM_3A = 256'hF1FFFFFEA7FE3C03E3B76FFFFF3FFFFF8F0E000000000000000F2FFFFFE71FF9;
defparam sp_inst_12.INIT_RAM_3B = 256'h8000000000007E1FFFFFC0FFCFE3309FA1FFFFE7FFFFFFE1E000000000000001;
defparam sp_inst_12.INIT_RAM_3C = 256'h7FFFFFFE03839FE007E0002007C3FFFFF80FFFEFF85CDBF3C3F3FFFFFFE31E3F;
defparam sp_inst_12.INIT_RAM_3D = 256'h8F1E6FE0FBF8CFFFFFFFE070078007F00007007E7FFFFF01FFFFFC78CCC3FBCE;
defparam sp_inst_12.INIT_RAM_3E = 256'hF8FFFFF837FE77E9EFE0F39FCF7FFFDFFF0E0018003F8000F31FC7FFFFC13FFF;
defparam sp_inst_12.INIT_RAM_3F = 256'h0F0003783FFF871FFFFC7DFF9FFD7F03FF23F9FFBFFBFF61C001C001FC001FFF;

SP sp_inst_13 (
    .DO({sp_inst_13_dout_w[30:0],sp_inst_13_dout[14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[14]})
);

defparam sp_inst_13.READ_MODE = 1'b0;
defparam sp_inst_13.WRITE_MODE = 2'b00;
defparam sp_inst_13.BIT_WIDTH = 1;
defparam sp_inst_13.BLK_SEL = 3'b000;
defparam sp_inst_13.RESET_MODE = "SYNC";
defparam sp_inst_13.INIT_RAM_00 = 256'hFFFFFE00000000000007FFFFFFFFFFFFFFFFFFFFF800F8783C07FFFFC0000000;
defparam sp_inst_13.INIT_RAM_01 = 256'hFFF0020018707DFFFFE00000000000007FFFFFFFFFFFFFFFFFFFFFC01E0E0381;
defparam sp_inst_13.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFE000007C60F1FFFFF00000000000001FFFFFFFFFFFFFFFFFF;
defparam sp_inst_13.INIT_RAM_03 = 256'h00000033FFFFFFFFFFFFFFFFFFFFF001FFF8F1C07FFFF00000000000001FFFFF;
defparam sp_inst_13.INIT_RAM_04 = 256'h003FFFF80000007F8007FFFFFFFFFFFFFFFFFFFFFF41FFFF1F8007FFFF000000;
defparam sp_inst_13.INIT_RAM_05 = 256'hFFFFFFFFFE3FC01FFFFF8000000004007FFFFFFFFFFFFFFFFFFFFFF87FFFF3F8;
defparam sp_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFE3FE0FCFFFF8000000000007FFFFFFFFFFFFFFFFFF;
defparam sp_inst_13.INIT_RAM_07 = 256'h00000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE7FE1F8FFFFC00000000000FFFFFF;
defparam sp_inst_13.INIT_RAM_08 = 256'hFF07FFFFF8000E00003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFC73F3E07FFFF0000;
defparam sp_inst_13.INIT_RAM_09 = 256'hFFFFFFFFFE0E1FC1FFFFFF800F800043FFFFFFFFFFFFFFFFFFFFFFFFFFFFF861;
defparam sp_inst_13.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFC0C07F3F3FFFFC01C0000C1FFFFFFFFFFFFFFFFFFF;
defparam sp_inst_13.INIT_RAM_0B = 256'h0000003FFFFFFFFFFFFFFFFFFC7FFFFFFFFE1F07F783FFFFE020000001FFFFFF;
defparam sp_inst_13.INIT_RAM_0C = 256'hE1F838FFFFE007800007FFFFFFFFFFFFFFFE3F8FFFFFFFFFE3FC3FC07FFFFE00;
defparam sp_inst_13.INIT_RAM_0D = 256'h1FFFFFFFFFC7EE0F8707FFFF03E00000FFFFFFFFFFFFFFFF87C1FFFFFFFFFC7F;
defparam sp_inst_13.INIT_RAM_0E = 256'hFFA3FFFFFC0C41FF3FFFFFF87C00FC00FFFFF0F800001FFFFFFFFFDFFFFFF0E0;
defparam sp_inst_13.INIT_RAM_0F = 256'hE600007FFFFFFFE0FFFFFFC1883F87FFFFFF0F030FC03FFFFFFE000003FFFFFF;
defparam sp_inst_13.INIT_RAM_10 = 256'hF871F1F9FFFFFDE03C0FFFFFFFFE1FFFFFF81107F9FFFFFFE0E1E07F07FFFFFF;
defparam sp_inst_13.INIT_RAM_11 = 256'h0FFFFFFFFFE33E0F1FFC0FFFFFFC0003FFFFFFFFC3FFFFFF00007FFFFFFFFF1C;
defparam sp_inst_13.INIT_RAM_12 = 256'hFF0BBFFFFE0001FFFFC3FFFC6603FBFE00FFBFFFC000FFFFFFFFF87FFFFFE000;
defparam sp_inst_13.INIT_RAM_13 = 256'hFF003FFFFFF9FE3177FFFFC0003FFF003FFF9E00FFEFE03FFFFFF8001FFFFFFF;
defparam sp_inst_13.INIT_RAM_14 = 256'h01FFE3F1FFFFFF8003FFFFFE0FC01FFFFFF00007FFC007FFF3C07FFEFE0FBFFF;
defparam sp_inst_13.INIT_RAM_15 = 256'h1FE003FFFFCE0018FF3F8FFFFBC0007FFFFFC1F003FFFFF600007FC001FFFE70;
defparam sp_inst_13.INIT_RAM_16 = 256'h800FFFFF800043F000FFFFF880010FFDFCFEFFF8003FFFFFF81E007FFFFCC000;
defparam sp_inst_13.INIT_RAM_17 = 256'h03FFFFFFFFE000017FFFF0001C38023FFFFFB0003997CFFFC7FE001FFFFFFF01;
defparam sp_inst_13.INIT_RAM_18 = 256'h00000FE3F0001FFFFFFFFFFE00002FFFFE003F000FE7FFFFE7E003007CFE7020;
defparam sp_inst_13.INIT_RAM_19 = 256'h03E31FEFFF9E000001FE3F001FFFFFFFFFFFC00000EFFFC01FE007C8FFFFFCF8;
defparam sp_inst_13.INIT_RAM_1A = 256'h00031FFE01FE03E04FF1FFF1C0000383F1F00FFFFFFFFFFFFC000018FFF007F8;
defparam sp_inst_13.INIT_RAM_1B = 256'hFFFFFFEFFFF8000023FF807E21F011FC1FFF7800000C7F9F81FFFFFFFFFFFF80;
defparam sp_inst_13.INIT_RAM_1C = 256'h000018FFE7FFFFFFF9E03FFC0000003FF80F0EF8067F007FCFE000018FF9FFBF;
defparam sp_inst_13.INIT_RAM_1D = 256'h0023F001FF18C0000003FF7FFFFFFF3803FF80000001FF0301FC009F800FF9EC;
defparam sp_inst_13.INIT_RAM_1E = 256'h000003C000078008FC003FE7000000007FF1FFFFFFFF8004F80000003E80203E;
defparam sp_inst_13.INIT_RAM_1F = 256'hFFFFFFC00000000000780000E0073F0007F8F00000000F7F9FFFFFFFFC000000;
defparam sp_inst_13.INIT_RAM_20 = 256'h0000000FFFFFFFFFFFFC7F4000000000000018018FC000FE1E58000003FFFCFF;
defparam sp_inst_13.INIT_RAM_21 = 256'h30F80001FC62000000007FFFFFFFFFFFEEFFE00000000004020063F0000FE3F8;
defparam sp_inst_13.INIT_RAM_22 = 256'h00000000000C3C3E00007F9C0000000007FFFFFFFFFFFE603FE0000000000040;
defparam sp_inst_13.INIT_RAM_23 = 256'hFFFFFFFE1800200000000001FC1FC0000FF1F0000000001FFFFFFFFFFFE3801F;
defparam sp_inst_13.INIT_RAM_24 = 256'h100000018FFFFFFFFFFFF0C0020000000000200FC00003FE3E0000000001FFFF;
defparam sp_inst_13.INIT_RAM_25 = 256'hFC71003FF8F00000000030FFFFFFFFFE3F078060000000000007F000007FC7C0;
defparam sp_inst_13.INIT_RAM_26 = 256'h000000000003FF2FE20FFF8FE009C080060FFFFFFFFF81F03FFC00000000000F;
defparam sp_inst_13.INIT_RAM_27 = 256'hFFFE1E003E000000000000003FFFF803FFF1FF0F00F00001EFFFFFFBE00FC038;
defparam sp_inst_13.INIT_RAM_28 = 256'hFFFC0000003FFFFFC3E000F000000000000007FFFE007FFE1FFFC3F8000005FF;
defparam sp_inst_13.INIT_RAM_29 = 256'hFFF007F1F8FFFFFC00003F1FFFFFF807E00FFE000000000000FFF7801F9FC3EF;
defparam sp_inst_13.INIT_RAM_2A = 256'h000000000003FFDE1FF87F1EFFFE00000FE7FFFFFFDC0041FFC000000000001F;
defparam sp_inst_13.INIT_RAM_2B = 256'hFFFF3F07FFFF0000000000007FF9C3FC03C3DFFC000001FDFFFFFFF3C01BFFF8;
defparam sp_inst_13.INIT_RAM_2C = 256'h0000000604FFFFFFFFF9FFE7F180000000001FFC7060000870700000003FFFFF;
defparam sp_inst_13.INIT_RAM_2D = 256'h1E000000000C00000001009FFFFFFFFFFFFC7E300003100003FC380000000838;
defparam sp_inst_13.INIT_RAM_2E = 256'h80060200001FF3C000000001000000066043FFFFFFFFFFFF9FCE001C3200007F;
defparam sp_inst_13.INIT_RAM_2F = 256'hFFFFFFFFFFCFC00000000007FFF0000000184000000082387FFFFFFFFFFFFEFD;
defparam sp_inst_13.INIT_RAM_30 = 256'h00000000F3FFFFFFFFFFFFFFF800000000007FEDE00001061180000000079FFF;
defparam sp_inst_13.INIT_RAM_31 = 256'h1800000000C0000000800C7FFFFFFFFFFFFFFF80000000000FF0E40000010620;
defparam sp_inst_13.INIT_RAM_32 = 256'h000000000E3F80000000003000000004400FFFFFFFFFFFFFFFF80000000021FC;
defparam sp_inst_13.INIT_RAM_33 = 256'hFFFFFFFFFFE38000000001C0FE00000000FC000000000000FFFFFFFFFFFFFFFE;
defparam sp_inst_13.INIT_RAM_34 = 256'h000000000CFFFFFFFFFFFFF07C00000000301F800000003FC000000000107FFF;
defparam sp_inst_13.INIT_RAM_35 = 256'h00000006FC0000000003800FFFFFFFFFFFFC3F800000000606700000001FF000;
defparam sp_inst_13.INIT_RAM_36 = 256'h00000000300080000600FF000000000270F0FFFFFFFFFFFFFFF000000001804E;
defparam sp_inst_13.INIT_RAM_37 = 256'hFFFFFFFFFFFF800000000E00000003801FC000000000E61E0FFFFFFFFFFFFFFE;
defparam sp_inst_13.INIT_RAM_38 = 256'h000000FB001FFFFFFFFFFFFFE000000001C0000003E007F0000000000E5801FF;
defparam sp_inst_13.INIT_RAM_39 = 256'h00F003EE00000000000FC701FFFFFFFFFFFF7F000000003C0F0001F007F80000;
defparam sp_inst_13.INIT_RAM_3A = 256'h00000000A000000003F780000000000070E1FFFFFFFFFFFFFFF0200000070000;
defparam sp_inst_13.INIT_RAM_3B = 256'hFFFFFFFFFFFF8000000000000000C0FFC00000000000001C1FFFFFFFFFFFFFFE;
defparam sp_inst_13.INIT_RAM_3C = 256'h00000001F07FFFFFF81FFFDFF800000000000000007CE00C00000000001C81FF;
defparam sp_inst_13.INIT_RAM_3D = 256'h701E701F0000000000001E0FFFFFF80FFFF8FF800000000000000078F03C0000;
defparam sp_inst_13.INIT_RAM_3E = 256'h000000003000080FF01F00000000002000C1FFFFFFC07FFF0CE0000000010000;
defparam sp_inst_13.INIT_RAM_3F = 256'hFFFFFC07C000780000007C00000180FC00000000000400983FFFFFFE03FFE000;

SP sp_inst_14 (
    .DO({sp_inst_14_dout_w[30:0],sp_inst_14_dout[15]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,ad[14]}),
    .AD(ad[13:0]),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15]})
);

defparam sp_inst_14.READ_MODE = 1'b0;
defparam sp_inst_14.WRITE_MODE = 2'b00;
defparam sp_inst_14.BIT_WIDTH = 1;
defparam sp_inst_14.BLK_SEL = 3'b000;
defparam sp_inst_14.RESET_MODE = "SYNC";
defparam sp_inst_14.INIT_RAM_00 = 256'h0000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0787C000000000000000;
defparam sp_inst_14.INIT_RAM_01 = 256'hFFFFFDFFFF8000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1F1FC00;
defparam sp_inst_14.INIT_RAM_02 = 256'hFFFFFFFFFFFFFFFFFFFFFFF8000000000000007FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000FFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_04 = 256'h0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE000000000000001;
defparam sp_inst_14.INIT_RAM_05 = 256'hFFFFFFFFFFC000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sp_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFFFFFFC00000000000000FFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000001FFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_08 = 256'h00000000000071FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF800000000000003;
defparam sp_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sp_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000000003FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000001FFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_0C = 256'h000000000000F87FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000007;
defparam sp_inst_14.INIT_RAM_0D = 256'hFFFFFFFFFFF80000000000001C1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sp_inst_14.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFFFFFFFFFFF8000000000000307FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_0F = 256'h19FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000001FFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_10 = 256'h000000000000021FC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000;
defparam sp_inst_14.INIT_RAM_11 = 256'hFFFFFFFFFFFC0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0;
defparam sp_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFFFFFFFFF80000000000000003FFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_13 = 256'h00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE00000000000000007FFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_14 = 256'h000000000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00000000000000;
defparam sp_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFF0000000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF80;
defparam sp_inst_14.INIT_RAM_16 = 256'hFFFFFFFFFFFFBFFFFFFFFFFF0000000000000007FFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFE3FFFDFFFFFFC000000000000001FFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_18 = 256'h000000000007FFFFFFFFFFFFFFFFFFFFFFFFC0FFF01FFFFFF80000000000001F;
defparam sp_inst_14.INIT_RAM_19 = 256'hFC00FFFFFFE0000000000000FFFFFFFFFFFFFFFFFFFFFFFFE01FF807FFFFFF00;
defparam sp_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFE01FC003FFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFF807;
defparam sp_inst_14.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFF81DE000FFFFFFF80000000000003FFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_1C = 256'h00000000000FFFFFFFFFFFFFFFFFFFFFFFF0F10001FFFFFFF00000000000007F;
defparam sp_inst_14.INIT_RAM_1D = 256'h001FFFFFFFE0000000000001FFFFFFFFFFFFFFFFFFFFFFFCFE00007FFFFFFE00;
defparam sp_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFFF80007FFFFFFF80000000000003FFFFFFFFFFFFFFFFFFFFFFFDFC0;
defparam sp_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFF0000FFFFFFFF00000000000007FFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_20 = 256'h00000000001FFFFFFFFF80BFFFFFFFFFFFFFE0007FFFFFFFE0000000000000FF;
defparam sp_inst_14.INIT_RAM_21 = 256'h0FFFFFFFFF80000000000003FFFFFFFFF0001FFFFFFFFFFBFC001FFFFFFFFC00;
defparam sp_inst_14.INIT_RAM_22 = 256'hFFFFFFFFFFF003FFFFFFFFE00000000000007FFFFFFFFF80001FFFFFFFFFFF80;
defparam sp_inst_14.INIT_RAM_23 = 256'hFFFFFFFFE0001FFFFFFFFFFE03FFFFFFFFFE0000000000000FFFFFFFFFFC0000;
defparam sp_inst_14.INIT_RAM_24 = 256'h00000000003FFFFFFFFFFF0001FFFFFFFFFFDFFFFFFFFFFFC0000000000001FF;
defparam sp_inst_14.INIT_RAM_25 = 256'hFFFFFFFFFF00000000000007FFFFFFFFFFF8001FFFFFFFFFFFFFFFFFFFFFF800;
defparam sp_inst_14.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFFF0000000000000FFFFFFFFFFFFC003FFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_27 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000001FFFFFFFFFFFFFC7;
defparam sp_inst_14.INIT_RAM_28 = 256'h00000000007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0000000000003FF;
defparam sp_inst_14.INIT_RAM_29 = 256'hFFFFFFFFFF0000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC00;
defparam sp_inst_14.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFFE1000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_2B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC2000000000003FFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_2C = 256'h0000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8F800000000007FF;
defparam sp_inst_14.INIT_RAM_2D = 256'hFFFFFFFFFFF000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7C0;
defparam sp_inst_14.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFFE000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_2F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE78000000000007FFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_30 = 256'h0000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9E000000000000FFF;
defparam sp_inst_14.INIT_RAM_31 = 256'hFFFFFFFFFF0000000000003FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF800;
defparam sp_inst_14.INIT_RAM_32 = 256'hFFFFFFFFF1FFFFFFFFFFFFC0000000000007FFFFFFFFFFFFFFFFFFFFFFFFDFFF;
defparam sp_inst_14.INIT_RAM_33 = 256'hFFFFFFFFFFFFFFFFFFFFFE3FFFFFFFFFFF00000000000000FFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_34 = 256'h0000000003FFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFFFFFFC00000000000001FFF;
defparam sp_inst_14.INIT_RAM_35 = 256'hFFFFFFF9000000000000007FFFFFFFFFFFFFFFFFFFFFFFF9FFFFFFFFFFE00000;
defparam sp_inst_14.INIT_RAM_36 = 256'hFFFFFFFFCFFFFFFFF9FF000000000000000FFFFFFFFFFFFFFFFFFFFFFFFE7FFF;
defparam sp_inst_14.INIT_RAM_37 = 256'hFFFFFFFFFFFFFFFFFFFFF1FFFFFFFC7FE000000000000001FFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_38 = 256'h0000000007FFFFFFFFFFFFFFFFFFFFFFFE3FFFFFFC1FF8000000000000003FFF;
defparam sp_inst_14.INIT_RAM_39 = 256'hFF0FFC1000000000000000FFFFFFFFFFFFFFFFFFFFFFFFC3FFFFFE0FF8000000;
defparam sp_inst_14.INIT_RAM_3A = 256'hFFFFFFFF5FFFFFFFFC08000000000000001FFFFFFFFFFFFFFFFFDFFFFFF8FFFF;
defparam sp_inst_14.INIT_RAM_3B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000000000000003FFFFFFFFFFFFFFFF;
defparam sp_inst_14.INIT_RAM_3C = 256'h000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8300000000000000007FFF;
defparam sp_inst_14.INIT_RAM_3D = 256'hFFE1800000000000000001FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF8700000000;
defparam sp_inst_14.INIT_RAM_3E = 256'hFFFFFFFFCFFFFFF00000000000000000003FFFFFFFFFFFFFFFFFFFFFFFFEFFFF;
defparam sp_inst_14.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFF83FFFFFE00000000000000000007FFFFFFFFFFFFFFFF;

SP sp_inst_15 (
    .DO({sp_inst_15_dout_w[29:0],sp_inst_15_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_15.READ_MODE = 1'b0;
defparam sp_inst_15.WRITE_MODE = 2'b00;
defparam sp_inst_15.BIT_WIDTH = 2;
defparam sp_inst_15.BLK_SEL = 3'b010;
defparam sp_inst_15.RESET_MODE = "SYNC";
defparam sp_inst_15.INIT_RAM_00 = 256'h12AC843A3AB2FE5468D3149014F0FFCFC0554505001646AC7C0EF5C56C5BC055;
defparam sp_inst_15.INIT_RAM_01 = 256'h14415545BFB0EB5705B1AAF1556B054EAB1504B8852900D0702FB951B00F3FFE;
defparam sp_inst_15.INIT_RAM_02 = 256'h30153900EAF1BED62B16ABBD5DE51BB0E8AC6F938A2705461B100FAC3F000554;
defparam sp_inst_15.INIT_RAM_03 = 256'h3B912FB74CB040FAF00300C6A451555A41A9B3F14F0AC55AC15AFF1AA41690BD;
defparam sp_inst_15.INIT_RAM_04 = 256'hB5F0316BC16C16AAAB0EFF8F556EA5380030CB0C422B1F14529E9508039EC6F9;
defparam sp_inst_15.INIT_RAM_05 = 256'h5AFD06DABAA4E6A45E4E9155539BFD24E406FC03FC00000F1A46AAAAA955A95B;
defparam sp_inst_15.INIT_RAM_06 = 256'h03FC0014F0645AEAD66FE555ABC303186C1BC0000FA4E869814E3A9534FAC060;
defparam sp_inst_15.INIT_RAM_07 = 256'h55514006FF9355B05534EBC2068413C6B0503EAE3A1D4FABEAAB8E4890F1ABFF;
defparam sp_inst_15.INIT_RAM_08 = 256'hE262B4FEBE56A984255F1BFFFC03FC004FC1419BAF95BCE91BAE0CFA5015AF00;
defparam sp_inst_15.INIT_RAM_09 = 256'h96AB456CE96EA7DEB53A56ABFC5AABF0005A9314EC55393F086ABE8F156B3F9B;
defparam sp_inst_15.INIT_RAM_0A = 256'h54F0000E431DFF683C501AA5591183DEABE4C0893A5A41BFFFFC03FC55301405;
defparam sp_inst_15.INIT_RAM_0B = 256'hB53F006FFEBFF15301A0143C519A5EA5BEBF9BE51A815AA56AEBC5555003015B;
defparam sp_inst_15.INIT_RAM_0C = 256'hA56A16BFEAABFFC195000FFAAB1AC0F002518AC308A000114049CFAE7AA9F049;
defparam sp_inst_15.INIT_RAM_0D = 256'h0EA05BC04FFF8CF5A5FE7AD4D1D05517FFC3FFF14C554404F295696AAABACE6F;
defparam sp_inst_15.INIT_RAM_0E = 256'hC031501413DA55A55BBEABFA5AAA95AFC0FFFC0005BA554FE50022C0F043EACB;
defparam sp_inst_15.INIT_RAM_0F = 256'h0016FEA943E94FE2C3F0043BCBF965D6FCE6A8B21E40F8B14DDD3C55BFFF00FF;
defparam sp_inst_15.INIT_RAM_10 = 256'hD0A90E95B88863C6B1FFFAC30FFF0450540C555A915AFA96A9697A5AFFC00000;
defparam sp_inst_15.INIT_RAM_11 = 256'h5545AAA5AABF9973ABFFFC0054555ABEE9543E4076FFFC003F06F9BC51BE569C;
defparam sp_inst_15.INIT_RAM_12 = 256'h38B1B0FABFF01C0D0025A4154DFA93F9AF88891B0607FFFC3FFFFC5540541541;
defparam sp_inst_15.INIT_RAM_13 = 256'h7C701AAAFFAFFFF04000055955001AEA5639BE64CEAFFFABC154555556FFFA5E;
defparam sp_inst_15.INIT_RAM_14 = 256'h91BABFFEAABC00005002AFFF9395A1B3905BCF6F39C366835561143AAA94D87A;
defparam sp_inst_15.INIT_RAM_15 = 256'h6BE5F8293C5B6C4FFAA8E9DC6B33141AABFABFFFC0004F15A55431AFA56C25A6;
defparam sp_inst_15.INIT_RAM_16 = 256'h003F55431A91550AA90AC3990AA55BFFFA96AF00F000015BFE953F06CE401AFD;
defparam sp_inst_15.INIT_RAM_17 = 256'hFFF055415540055A6F3F96A6C546F9AAE4F5B84000FFB552373B71546AAFAAFC;
defparam sp_inst_15.INIT_RAM_18 = 256'h40FFF924213C226A56AAAAAFFF03F154005A95A57A558EA9642FF9AFFEBAAAAF;
defparam sp_inst_15.INIT_RAM_19 = 256'h56A5560FA6A57FE9FF0FEAAAFFFFF00405540003FFC56B00EAAB06C8964FD660;
defparam sp_inst_15.INIT_RAM_1A = 256'h3FFAAC6154396BDAE716E913F4FFAA4F9E1D2C16A96A59AFFFFFFF1540551941;
defparam sp_inst_15.INIT_RAM_1B = 256'hBFAAA966BFFFFF305501A400C06956983FAAA47F97FF0FAAAAAAABFF00055014;
defparam sp_inst_15.INIT_RAM_1C = 256'h756FCFFE9595555AAB00000000FFF95DC050FF3F014E1B823E0EA94E5521D3F5;
defparam sp_inst_15.INIT_RAM_1D = 256'h00F0392DED38E54E903A623FF3BFFEF99BBFFEB000151553F01568165AA2B950;
defparam sp_inst_15.INIT_RAM_1E = 256'hF300506500C1B956FA45B6F95686FF3FAAA554500596AFAF0FCFCFA472FEFF10;
defparam sp_inst_15.INIT_RAM_1F = 256'h001555556ABFFFFFA562901B0FFFCF84891B85C094FE5377AFCDAFABEAAFFFFF;
defparam sp_inst_15.INIT_RAM_20 = 256'hBD3E550E226C856AABEAB03F3FFFC00195100B3A58D50B98F4A91ABFFFFEA550;
defparam sp_inst_15.INIT_RAM_21 = 256'hFD2E456EB3E7FAA6BFFFFFA50000569555556AA9AA5440FF0696FFA4FE3EB1BE;
defparam sp_inst_15.INIT_RAM_22 = 256'h55654626AC00F2E54FE40F51695350154DED635555AFAAC030FFFFC00555417F;
defparam sp_inst_15.INIT_RAM_23 = 256'h955AAA96C0003C003F145A56AAAAF65A6FFFFC00DAFFFFAAA500016AA5554001;
defparam sp_inst_15.INIT_RAM_24 = 256'h0F3FFFFA5AA55006AAF9554000015535C32F0FFCF0339FEC0003940069389D7D;
defparam sp_inst_15.INIT_RAM_25 = 256'hABFFB93929BE5500156BE203F66A6BAAAAF00001543050696AA56B99BEBEC0FC;
defparam sp_inst_15.INIT_RAM_26 = 256'h0040059555A5AABFAACF2B17FEACBFFFFAAAAA5006AAAA550C3C30573FF70ABE;
defparam sp_inst_15.INIT_RAM_27 = 256'h541AAAAA943FFFF0B37FFFB00016554E524153C155AA994941DAA9AAABEAF001;
defparam sp_inst_15.INIT_RAM_28 = 256'h1BFFF9D0F91C6AAAAAAFAAC00530F3C6550156FAC3AB00FC5FE5BEFFF0FEABFE;
defparam sp_inst_15.INIT_RAM_29 = 256'hB980973C0FAFEBEF00C3FFFFFEA56AAAAA54FFF0C6353D58555BFEAE903C0553;
defparam sp_inst_15.INIT_RAM_2A = 256'hC01A44F6B4FFDA91A00C1ABFFA805F9E43E57155AAAAAFFFF054FEFC154001AA;
defparam sp_inst_15.INIT_RAM_2B = 256'h56AAAFFFFEF1500C0F15551556FABEAFAFFAD3EB3C50FFFFFCFFE9AAAAA950FF;
defparam sp_inst_15.INIT_RAM_2C = 256'hACF00FAAFC000FAAAAAAA5503BC05FCFCA793F1AAA955625A59050392540FB05;
defparam sp_inst_15.INIT_RAM_2D = 256'h8054F0C63C3FE54393955A955556AABFFFFFC555553F1056A5AAEB9BF97C3F3F;
defparam sp_inst_15.INIT_RAM_2E = 256'h95503F002A9BBE725AE5853EACEFF03FABF000FAAAA5655554FF051BFAEA524C;
defparam sp_inst_15.INIT_RAM_2F = 256'hAAAA9555565030126FEB7F34D36F3EAAB10403A53A3AAAC579655AAABFCF3F55;
defparam sp_inst_15.INIT_RAM_30 = 256'h9394EFF1C47AA96AAAFFFC055155453F04A96AB3F95B0984EE640AFFFEABC00E;
defparam sp_inst_15.INIT_RAM_31 = 256'hFCE47CE6F07FFAEBAF3FFFF03E941A55555554005FC3A1C14E3DC54000555503;
defparam sp_inst_15.INIT_RAM_32 = 256'h15414E871A439769569554000E4D3FFC61F87EA6AAABFFFC150140040306A6F6;
defparam sp_inst_15.INIT_RAM_33 = 256'hAAAEBFFFF0540003C1401A9BEAB0E5C3ECB5035AFFFCFFFFFC3E955555555A95;
defparam sp_inst_15.INIT_RAM_34 = 256'hB00FFFFFFFFFFEA555AA5A6A9555550F1CAA53AD502A9543FFF4D3ABF76C363A;
defparam sp_inst_15.INIT_RAM_35 = 256'hFCEB55553FAB9D3FF0B7002D3EBABFFFFFC0450003C665A5199180EB00FF0009;
defparam sp_inst_15.INIT_RAM_36 = 256'h500306AA955A45BFF033E83CEAAFFEA6BFFFFEAAA956BFB9559555550C21AA5F;
defparam sp_inst_15.INIT_RAM_37 = 256'hAFAAAAFFE95696956540B1BA4FE4F71410E8C5E3FC6D8553B43FFAFFFCFAF105;
defparam sp_inst_15.INIT_RAM_38 = 256'h0FCB61AA93D0FFEBFFFFFFC40540545AAA59591AFC3FF030ABFE6BAA96ABFFFE;
defparam sp_inst_15.INIT_RAM_39 = 256'h6B00AAC103ECFD6AAAAAABFFFEFEFAAAFA95595555A545B1AA438E82FFE9086E;
defparam sp_inst_15.INIT_RAM_3A = 256'h45569556B0154E400641FF7B10C1871BFF92D3FFFFFFFFCFC0C5016566A6A565;
defparam sp_inst_15.INIT_RAM_3B = 256'hFFFABCFF0FF30406A81B9AAAFA58CEAB0FC403F9AAAAAAAAAFFFFBFFEAA95555;
defparam sp_inst_15.INIT_RAM_3C = 256'hA5AAAAAAAAAFFFFFFFEA955555016A555AABC640FAA4E9575BC06DB1AC0F9180;
defparam sp_inst_15.INIT_RAM_3D = 256'h5500E93A9EBF162DAABC0F8B40FFFBFFFCFBC05415957395656A771FECFBFD43;
defparam sp_inst_15.INIT_RAM_3E = 256'h500541FF9555AF0F303F9FB0FE954055566AAFFFFFFFA95505640569555A96DA;
defparam sp_inst_15.INIT_RAM_3F = 256'hABFEFE955506A95AA555AA46D550143FAA7FAAB2DBFBFC0E2D50FFFFFFFFEB04;

SP sp_inst_16 (
    .DO({sp_inst_16_dout_w[29:0],sp_inst_16_dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_16.READ_MODE = 1'b0;
defparam sp_inst_16.WRITE_MODE = 2'b00;
defparam sp_inst_16.BIT_WIDTH = 2;
defparam sp_inst_16.BLK_SEL = 3'b010;
defparam sp_inst_16.RESET_MODE = "SYNC";
defparam sp_inst_16.INIT_RAM_00 = 256'h3EAB8695400555553A6F00FFFFAFAABABFFFFFFFFFFFFFFC3C0FF0C0FC001555;
defparam sp_inst_16.INIT_RAM_01 = 256'hFFFFFFFFFFF0FF0303F000055555AAA555AAAA416A9555000555400005504000;
defparam sp_inst_16.INIT_RAM_02 = 256'h9AAA9555000555003F0000000FAAAA1A550155540EAF000EAAFFFAABEAFFFFFF;
defparam sp_inst_16.INIT_RAM_03 = 256'h43FF003EA6AFFFAAAFFEFFBFFFFFFFFFFFFFF3F00F0FC000155555AAAAAAAAAA;
defparam sp_inst_16.INIT_RAM_04 = 256'hF0F030001556AAAAAAFAAAA5AAAAAA95554515A503EAFF0003FAAAADA9501555;
defparam sp_inst_16.INIT_RAM_05 = 256'hA4FAAABFFFFFAAAA86A555555400003FAAAAABFEABFFFFFAFFFFFFFFFFFFFFFF;
defparam sp_inst_16.INIT_RAM_06 = 256'hFEABFFFFAFFFFFFFFFFFFFFFFFC3030156AABFFFFAAA56AA55505AAA9500155A;
defparam sp_inst_16.INIT_RAM_07 = 256'hAAAAAAAAAAA9555AAA950015AAA4E96AAFFFEAAA966AA5555555500FAA5AAAAA;
defparam sp_inst_16.INIT_RAM_08 = 256'hA95DAA555555550FEAA5AAAAABFEABFFFABFFFFFFFFFFCFFFFFF0CFD555555AA;
defparam sp_inst_16.INIT_RAM_09 = 256'hFFFFFFFCFFFFFFFFF54000000155555AAAAAA9AA56AA954056AA93A5AAAAEAAA;
defparam sp_inst_16.INIT_RAM_0A = 256'hAA5AAAA55456AA9396AAAAAAAA958AA55555150FEAAAAAAAAAABFEABFFEFFFFF;
defparam sp_inst_16.INIT_RAM_0B = 256'hEA95AAAAAAAAAFFEFFFFFFEBFFFFFFFFFFFFFFFFFFC000000000155555545555;
defparam sp_inst_16.INIT_RAM_0C = 256'hFFFF0000000000155555500000556A5AA9556ABE9E5AAAAAAAA5176A95550550;
defparam sp_inst_16.INIT_RAM_0D = 256'hFA4E556AA5555176AA55401503AAAAAAAABEAAAFFBFFFFFFAFFFFFFFFFFFCFFF;
defparam sp_inst_16.INIT_RAM_0E = 256'hBFEFFFFFFEBFFFFFFFFFFFFFFFFFFC0015000155555555500000056A5AA9556A;
defparam sp_inst_16.INIT_RAM_0F = 256'h5555555554000FC5695AAA956AAA4E555655550B6AAA550550FA96AAAAAAFFAA;
defparam sp_inst_16.INIT_RAM_10 = 256'h76AAA555550F94155AAAAABEFAAAFFFFFFFBFFFFFFFFFFFFFFFFFFF000155555;
defparam sp_inst_16.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFF3C00001555555555555554000055556AA95AAAA4F95555551;
defparam sp_inst_16.INIT_RAM_12 = 256'h3C055A55555AABFA93955555571AA9555550FA9055AAAAABEAAAABFFFFFFFFFF;
defparam sp_inst_16.INIT_RAM_13 = 256'h415AAAAAAAAAAAAFFFFFFFFFFFFFFFFFFF3FFFFFCF0000001555555555555550;
defparam sp_inst_16.INIT_RAM_14 = 256'hFFFC0000000155555555555554000559555565AAEA5295545561AA9555550F95;
defparam sp_inst_16.INIT_RAM_15 = 256'hAAAA4F954155C6A5555500FA4045AAAAAAAAAAAABFFFFAFFFFFFEFFFFFFC3FFF;
defparam sp_inst_16.INIT_RAM_16 = 256'hFFEAFFFEFFFFFFFFFFFFC3FFFFFFF00000000055055555555555405565555556;
defparam sp_inst_16.INIT_RAM_17 = 256'h0005555555555555559555556AAAAA4E5505586AAA554003E9405AAAAAAAAAAB;
defparam sp_inst_16.INIT_RAM_18 = 256'hAA5555403E9695AAAAAAAAAAAAFEAFFFFFFFFFFFFFFFCFFFFFFFFFC000000000;
defparam sp_inst_16.INIT_RAM_19 = 256'hFFFFFF0FFFFFFFFF005000000000055555555554001555AA5555AABA4E5015B6;
defparam sp_inst_16.INIT_RAM_1A = 256'h4000015AAA95556AA94E55AF1A5555500FE556AAAAAAAAAAAAAAAAFFFFFFFFFF;
defparam sp_inst_16.INIT_RAM_1B = 256'hAAAAAAAAAAAAAAEFFFFFFFFFBFFFFFFC3FFFFFFFFC0050000000000055555555;
defparam sp_inst_16.INIT_RAM_1C = 256'hFFF010000000000000555555550000016AAA5595AAA54EAAF1A55550003E5406;
defparam sp_inst_16.INIT_RAM_1D = 256'hAA5A954FAB065550003FE94005AAAAAAAAAAAAAFFFFFFFFEAFFFFFFFFFF3FFFF;
defparam sp_inst_16.INIT_RAM_1E = 256'hAEFFFFFFFFBFFFFFFFFFFFFFFFFFC040000000000000000050101000055555AA;
defparam sp_inst_16.INIT_RAM_1F = 256'h000000000000000000055555A55565550FFF151500FFFE940016AAAAAAAAAAAA;
defparam sp_inst_16.INIT_RAM_20 = 256'h003FFFFA94016AAAAAAAAFEAEAAABFFFFFFFFF3FFCFFFFFCFFFFFF0000000000;
defparam sp_inst_16.INIT_RAM_21 = 256'hFFFFFFFFF3FFFFFC0000000000000000000000000000150055555555003FF000;
defparam sp_inst_16.INIT_RAM_22 = 256'h000000400155055550000F000003FFFFFA5005AAAAAAAABFEFAAAABFFFFFFFFF;
defparam sp_inst_16.INIT_RAM_23 = 256'hAAAAAAAABFFFEBFFEAFFFFFFFFFFFFFFFFFFFC00F00000000000000000000000;
defparam sp_inst_16.INIT_RAM_24 = 256'h0F000000000000000000000000000004C300500105440FFC0003FFFFFFEA5006;
defparam sp_inst_16.INIT_RAM_25 = 256'h0000003FFFFFFFFFFFFEA9541AAAAAAAAAAFFFFFFFEFFFFFFFFFFFFFFFFFC0FC;
defparam sp_inst_16.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFCF3F03FFFC000000000000000000000C3C30004FFF0000;
defparam sp_inst_16.INIT_RAM_27 = 256'h00000000003FFFF0043FFFF00000000FFEFFFEBFFFFFFAA5556AAAAAAAAAAFFF;
defparam sp_inst_16.INIT_RAM_28 = 256'hFFFFFFAA5556AAAAAAAAAABFFFEFAEBFFFFFFFFFC3FF00FC0FFFFC0005000000;
defparam sp_inst_16.INIT_RAM_29 = 256'hFFC0FF3C0FFFFFF055140000000000000000FFF0C0403C0FFFFFFFFFFFEBFFFE;
defparam sp_inst_16.INIT_RAM_2A = 256'hC00000F03FAABFFFFFFBFFFFFFC00FFAA9555AAAAAAAAAAAAFFFAAABFFFFFFFF;
defparam sp_inst_16.INIT_RAM_2B = 256'hAAAAAAAAAAAFFFFBFAFFFFFFFFFFFFFFFFFFC3FF0155000001000000000000FF;
defparam sp_inst_16.INIT_RAM_2C = 256'hFC05500001555000000000003FC00FCFC03FEAFFFFFFFF000000003FEAAA55AA;
defparam sp_inst_16.INIT_RAM_2D = 256'hC000F0C041400003FEAAAAAAAAAAAAAAAAAABFFFFFEAFFFFFFFFFFFFFFFC3F3F;
defparam sp_inst_16.INIT_RAM_2E = 256'hFFFFEAFFFFFFFFF3FFFFC03FFCFC0540000555000000000000FF003FFFC003FB;
defparam sp_inst_16.INIT_RAM_2F = 256'h0000000000003003FFFF0040FF004000055554003FEAAABFEAAAAAAAAABAEAFF;
defparam sp_inst_16.INIT_RAM_30 = 256'h03FFAAAFC0EAAAAAAAAAABFFFFFFFFEAFFFFFFF3FFFF0FC0FFF0000000001550;
defparam sp_inst_16.INIT_RAM_31 = 256'hFCFFFCFFF03FFFC00040000540000000000000000FC3F015503C155555555554;
defparam sp_inst_16.INIT_RAM_32 = 256'h00000FC05554005555555555500FEAABF000EAAAAAAAAAABFFFFFFFFFEFFFFFF;
defparam sp_inst_16.INIT_RAM_33 = 256'hAAAAAAAAAFFFFFFEBFFFFFFFFFF0FFC3FCF003FF000100000140000000000000;
defparam sp_inst_16.INIT_RAM_34 = 256'hF150000000000000000000000000000F01555401555555540000FEAAAF0143EA;
defparam sp_inst_16.INIT_RAM_35 = 256'h0100555540000FEAAFF0554FEAAAAAAAAABFFFFFFEBFFFFFFFFFC0FF00FF000F;
defparam sp_inst_16.INIT_RAM_36 = 256'hFFFEFFFFFFFFFFFFF033FC3CFFF000000000000000000000000000000C055550;
defparam sp_inst_16.INIT_RAM_37 = 256'h0000000000000000000005555000F0555500C0FEABFC15543FEAAAAAABAAAFFF;
defparam sp_inst_16.INIT_RAM_38 = 256'hFABF055554FFAAAAAAAAAABFFFFFFFFFFFFFFFFFFC3FF030FFFFC00000000000;
defparam sp_inst_16.INIT_RAM_39 = 256'hFF00FFC003FCFF000000000000000000000000000000000555540FC000000FFF;
defparam sp_inst_16.INIT_RAM_3A = 256'h00000000055550000000FFEAFFBFC0555554FEAAAAAAAABABFBFFFFFFFFFFFFF;
defparam sp_inst_16.INIT_RAM_3B = 256'hAAAAABAAFAAEFFFFFFFFFFFFFFFCCFFF0FC003FC000000000000000000000000;
defparam sp_inst_16.INIT_RAM_3C = 256'hF0000000000000000000000000000000000015550000FFFEAABFFC0556A554FF;
defparam sp_inst_16.INIT_RAM_3D = 256'h5555003FFAAAFF015556A553FFAAAAAAABAABFFFFFFFF3FFFFFFF30FFCFFFC03;
defparam sp_inst_16.INIT_RAM_3E = 256'hFFFFFFFFFFFFFF0F303FFFF0FFC0000000000000000000000000000000000015;
defparam sp_inst_16.INIT_RAM_3F = 256'h00000000000000000000000015555540003FFFF0155556A54FFFAAAAAAAAAAFF;

SP sp_inst_17 (
    .DO({sp_inst_17_dout_w[29:0],sp_inst_17_dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]})
);

defparam sp_inst_17.READ_MODE = 1'b0;
defparam sp_inst_17.WRITE_MODE = 2'b00;
defparam sp_inst_17.BIT_WIDTH = 2;
defparam sp_inst_17.BLK_SEL = 3'b010;
defparam sp_inst_17.RESET_MODE = "SYNC";
defparam sp_inst_17.INIT_RAM_00 = 256'hEA0A3D7FDFDFFF7DC0A07D88882A00222A2A00208A20A081615227BF01F77D5F;
defparam sp_inst_17.INIT_RAM_01 = 256'h2200AA020A05AA7C5605D7DDF5D577D5DDFD55D7D75D5F5DD555F7D55D75D577;
defparam sp_inst_17.INIT_RAM_02 = 256'hDFDFD755F7777D55C87D57FFDA82AA55DFFDDF55F2A0DF708002A20A88080288;
defparam sp_inst_17.INIT_RAM_03 = 256'h5400F5C2202AA2208A28802820208AAA82208607DA5A1FF5F7F7FDD577D7DD55;
defparam sp_inst_17.INIT_RAM_04 = 256'h25874777D7DFDD555F5D5FDF75F55DF5DD775DDFDE82A2F756A8000375D7F7D5;
defparam sp_inst_17.INIT_RAM_05 = 256'h55820A82888A08A0B77D7777D7F555C808080808A8A28820AAA228A008A2A2A8;
defparam sp_inst_17.INIT_RAM_06 = 256'hA882A082228820A8202220A202BE56755D77775F57D7D5DDD5D755777F7F55DD;
defparam sp_inst_17.INIT_RAM_07 = 256'h7FD57FFDFDD7D5D777D557D5F75F028A020A228280F75FF7FFF7FFD0AAA0AA02;
defparam sp_inst_17.INIT_RAM_08 = 256'h28A3D7FDDDD557728A80A808222022AA8022A208A02A098288A859817FF77DFD;
defparam sp_inst_17.INIT_RAM_09 = 256'h000A02A98A0028A82777FF5F7DD7FF5FFFD5FDFF5F5DF5D5D777540222220808;
defparam sp_inst_17.INIT_RAM_0A = 256'h75757DD55DDD7FF4AA00AAAA88281F7757DFD55002008082808208A2AA8A2A88;
defparam sp_inst_17.INIT_RAM_0B = 256'h2AA082020AA2888822A22882A08008AA8A82AA82281DFFFFD77DD57FD7F55FDF;
defparam sp_inst_17.INIT_RAM_0C = 256'h2020DD7F77FD55F75F5577F5FD7FFD57F577DDD5F08A802088A0AA5FF7F5DD77;
defparam sp_inst_17.INIT_RAM_0D = 256'h5D722A02AAA00A2F5D5DFD5FDE228088AA80828002A8800802A0A8A02A8A1282;
defparam sp_inst_17.INIT_RAM_0E = 256'h2A82222AA0282AA2082A08A28800ABDDF5DF7D5FDDD77FD5DF577DDFF775DFF5;
defparam sp_inst_17.INIT_RAM_0F = 256'hFFF77DFDDD5DD23FFF7FD775F5FD7AAA002200A05FDD77F77F2A2A008AA22820;
defparam sp_inst_17.INIT_RAM_10 = 256'h2577DDDF7FD0082820282A828A000802A22282822288AA8822A88287DFD5555F;
defparam sp_inst_17.INIT_RAM_11 = 256'hAAA8AA2A0228AA0C977FFDFFFFD55FD775FDD5FFF7FF5DF57FD77550A02AA202;
defparam sp_inst_17.INIT_RAM_12 = 256'h43FFF5D7DFFF57FF762228AAAA57575D55FD02A0880080A2880A80A288A82882;
defparam sp_inst_17.INIT_RAM_13 = 256'h2000222A2880A808002A8280AA2A00022A40AA22BA7DFDF5DD57D575FD7FDD55;
defparam sp_inst_17.INIT_RAM_14 = 256'h882BF5575F5DFF577DF5F5FDFFD7D5F7DF7775D7D574A00200AFFF57F7F5F0A2;
defparam sp_inst_17.INIT_RAM_15 = 256'hF7DD50AA8A22BF7FDFFD75A28A08282AA8A800002880A080A2088A82028BCA22;
defparam sp_inst_17.INIT_RAM_16 = 256'hA808A8200AA2AA88AA8A1EA80A282F55FF555757FDF557DF57F7D575DF75D75F;
defparam sp_inst_17.INIT_RAM_17 = 256'h57DDFDF7F5DFF55F57F57D5DDF75F5DA80AA035D55DD7DF488A00820A820A2AA;
defparam sp_inst_17.INIT_RAM_18 = 256'h55D5D57742082A8828000A220AA8888808800800222238A002200AB5D7DD5FF7;
defparam sp_inst_17.INIT_RAM_19 = 256'hA2220078008A0A8AF5FDD5FF5F555D7D5F7DD57DFD77D5F5DF5F757758880A27;
defparam sp_inst_17.INIT_RAM_1A = 256'hDD5DFD7757FFF7DDFD582A88775D575DD8AA020AA008002A200080A08A8208A2;
defparam sp_inst_17.INIT_RAM_1B = 256'h8A2AA8008082A2A8802AAA822A8028AB48AA00082BFFFDD557555F57555FF555;
defparam sp_inst_17.INIT_RAM_1C = 256'h2087FFD77F7FF5755DF57F5FFF7FD5DD5DF57D57F7D77AA0057D757F754228A0;
defparam sp_inst_17.INIT_RAM_1D = 256'hF5D5755A285DDD5D7F48200A8A02200808808228202A2000822002202A8682A2;
defparam sp_inst_17.INIT_RAM_1E = 256'h0A80AA0802280A8A0A08A8AAA2AA97F5FF5F775D777F575DF555575F5F57F5D7;
defparam sp_inst_17.INIT_RAM_1F = 256'hF5DDD5557D7FFD7DDF7D755F57F5FD7DFA287F5D5D228AA8028880A0282002A0;
defparam sp_inst_17.INIT_RAM_20 = 256'h7D422888A0288A08202A80A2A000A800822A8060A1A020A18088AAD557FFDDDF;
defparam sp_inst_17.INIT_RAM_21 = 256'h000A0A022CA80209D55FDF5D7F5D5FD77D55FFF5D77FDD5777D557DFF5E2ADFD;
defparam sp_inst_17.INIT_RAM_22 = 256'h7F77D77D7DD755D55F5D50DD755E22882200000A80202028880A08AA20800220;
defparam sp_inst_17.INIT_RAM_23 = 256'hAA82AA28822A82088828882228A800A88882A9DDA755FFF55DF5FDD57D5FFFFF;
defparam sp_inst_17.INIT_RAM_24 = 256'h58DF557DF55F5DF755F7D57555D7577D14D777D777775A01775400A888208828;
defparam sp_inst_17.INIT_RAM_25 = 256'h55FDDF4A02002A0AA8002228A20008A0A22A8A2AA88200A82808A82028A01D89;
defparam sp_inst_17.INIT_RAM_26 = 256'h2082A8AA08AA80A288B2EA742201F5555D55FFD77D57D7DDD9696DFFF0A2F7FD;
defparam sp_inst_17.INIT_RAM_27 = 256'hF7DD7F57F76AAAAD574A2285F5F5FD7A2828AA8AA8A8A0A2220A802A02208A0A;
defparam sp_inst_17.INIT_RAM_28 = 256'h02AA8A2A082A8800002AAAA0828A2A020A08AA22BE2857A970A82B55557FFF55;
defparam sp_inst_17.INIT_RAM_29 = 256'h201DA069D08A02A57755FF55F77FD7FFD5D722A5B7FDE1508020A2A28288A80A;
defparam sp_inst_17.INIT_RAM_2A = 256'hBD77FD8F4A8002A0202208AA82BD522A28A8A8800A8220028A8A0A822A8A2208;
defparam sp_inst_17.INIT_RAM_2B = 256'h002A2008A2202820A02A0820022020A02A8A9620775DFFFD57F5F55F57555FA0;
defparam sp_inst_17.INIT_RAM_2C = 256'h09F7F7D5F7FFFDF555555D5F60B77238BF6A2A220AA0227555D7D5C022220228;
defparam sp_inst_17.INIT_RAM_2D = 256'h3FD5AF17D7DDFDDC028AAA08A020A28A002A000200AA00A02AA8080808094268;
defparam sp_inst_17.INIT_RAM_2E = 256'h8A22A0A8220A28240A8015482383F75F77DF7FDFFF5FDFD5D7025FEAA8175C28;
defparam sp_inst_17.INIT_RAM_2F = 256'hD57F7FF57FDD6D5482A075F7085DDFD5D75D5D57EAA02A8AAA00A20A28202280;
defparam sp_inst_17.INIT_RAM_30 = 256'hD422080A1722A00A2A208208020808808882280408A25A1D280775F75D575D77;
defparam sp_inst_17.INIT_RAM_31 = 256'h8320A1A0A7622015575FD55FF77575FFFFFFD7D7723E0D57FFC955DFFDD7FF5F;
defparam sp_inst_17.INIT_RAM_32 = 256'hF5F57895DF5555FDF5755D5F7FFA8AA20FF52280AAA80000822A8A2008822AA0;
defparam sp_inst_17.INIT_RAM_33 = 256'h8A82A00002A0A080A0002882028728360107DC80FF5D7FD557F7755FFF557575;
defparam sp_inst_17.INIT_RAM_34 = 256'h855F7D5F5D757F5D55D7F7D5FD7557507FD57F7F775D757DDD552A082275F422;
defparam sp_inst_17.INIT_RAM_35 = 256'hD7FF57555F7DF08A028D5570220A82028228800AA822A222A0A2352AD52057DA;
defparam sp_inst_17.INIT_RAM_36 = 256'h228002A8A2008202A5642BE10A0DFDF75FF57D555555D7D7FF7DD5F75BD7DDF7;
defparam sp_inst_17.INIT_RAM_37 = 256'h7FF7F757DFDFFDD5F7F77D7DDF5D07F7DD5717020A0B7FDDE2200A200A8A02A8;
defparam sp_inst_17.INIT_RAM_38 = 256'hAA227FD5FD08A82800AA200888AAA80208022A2083E8056D2088B57FD7D7575F;
defparam sp_inst_17.INIT_RAM_39 = 256'h0A5F0A9D740908DFFFFF57D57FFF7F57FDF57FDFD5F5D5F5D7757037F5F7D0A0;
defparam sp_inst_17.INIT_RAM_3A = 256'h755FF575DDF755755F550002280A9F5757F782A0AA02A0208A2882002000A822;
defparam sp_inst_17.INIT_RAM_3B = 256'h800A8AA8A20A8888880A828288A9908A5A37F6AB7FFDF555FF7F7D55D55755FD;
defparam sp_inst_17.INIT_RAM_3C = 256'h2DF57F7FF57D5577FD557D55755F77FD57FDD75DD75D2000A88AA9F5D7F7FFA2;
defparam sp_inst_17.INIT_RAM_3D = 256'h7DFDF7C882A288DFFF755DF6A0000A008A8A028008800C2A8A8A06D8010A83DE;
defparam sp_inst_17.INIT_RAM_3E = 256'hA282A200A222A2786F62A0A5A297DFFFF77D7D7D555DDFF5FDFFF577F5D7DDF7;
defparam sp_inst_17.INIT_RAM_3F = 256'hFF5FD7FFD5F75FFF5F55F7DFFFF7D75FF7CA008DD57FD55D702A00A20200A88A;

SP sp_inst_18 (
    .DO({sp_inst_18_dout_w[29:0],sp_inst_18_dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]})
);

defparam sp_inst_18.READ_MODE = 1'b0;
defparam sp_inst_18.WRITE_MODE = 2'b00;
defparam sp_inst_18.BIT_WIDTH = 2;
defparam sp_inst_18.BLK_SEL = 3'b010;
defparam sp_inst_18.RESET_MODE = "SYNC";
defparam sp_inst_18.INIT_RAM_00 = 256'h23FCC43A4FC6F9431B64A9E510FFFFFEFF000030CF05315B2BF9A0B01BC5ABFF;
defparam sp_inst_18.INIT_RAM_01 = 256'h030000006AAF9603C06C156BFFC15AA4CC155491D94FA54ADAB08EAAC1400002;
defparam sp_inst_18.INIT_RAM_02 = 256'h016A52AA405A032B4C5BFFFEA2395BB0F8F17F9375D16A9C5B13FEABFBFC0010;
defparam sp_inst_18.INIT_RAM_03 = 256'h374C85DB81BF03EABFFFC3F19041000500556EAC0AC5BC056FF0016FE96AA5BE;
defparam sp_inst_18.INIT_RAM_04 = 256'hA0AF2F056FC16BFFFF0F0F9F556FFA4E6A996C11974C6069A79FEA5803A31AF9;
defparam sp_inst_18.INIT_RAM_05 = 256'hAF06AB2FCFF93BE95D4FD5A95246A7493556FC0FABFFCC3FC531955555005406;
defparam sp_inst_18.INIT_RAM_06 = 256'hFFBFFFC3EF100696855A95005ABEFEF6C1AF045003F901BAE6534BEE89406A81;
defparam sp_inst_18.INIT_RAM_07 = 256'hAAAA955BFFA7AA85AE4E406B1A95B96B15A543C34EC94FAFE55524E1E506AAFF;
defparam sp_inst_18.INIT_RAM_08 = 256'h376164FFCF5557624AA41BFBEF3FEFFF0FF030565A406BA4C65AFBABEAAF0156;
defparam sp_inst_18.INIT_RAM_09 = 256'h55A6441BA46A929AAE940055ABC00055556F901401AA43556CAE8329AEF050FC;
defparam sp_inst_18.INIT_RAM_0A = 256'hA9055654E572FF6E96FAAFFABF618E8EFFE3C374D3FF96BFFFBF0FAF00FF03C1;
defparam sp_inst_18.INIT_RAM_0B = 256'h639555BFFAAEBC0FF05300FF01555A50696E469406BC00001596B03FFEAAAABC;
defparam sp_inst_18.INIT_RAM_0C = 256'h955AC15A9556AAAF0FFFE95501AF155554EADBC30EC6AAAAA6920E952AA9FC27;
defparam sp_inst_18.INIT_RAM_0D = 256'h0EE9EC699005DC2050FA3AC3488EBE6BFFC0FEB00F010000F145151A9565FD1A;
defparam sp_inst_18.INIT_RAM_0E = 256'hFFF00303C3C6405456A9A6A916AA5416AFAAABFABC143FFA53FEF71505950F1B;
defparam sp_inst_18.INIT_RAM_0F = 256'hFFF05500FA90F9B7140569401BF9AAEB567F0DC2050FE7A03788E6FABFFF00FF;
defparam sp_inst_18.INIT_RAM_10 = 256'h1354FA5067776EAC06FFEAC3CEFFC003033F14154016A552981569556ABFFFFF;
defparam sp_inst_18.INIT_RAM_11 = 256'h0031559069AA457F55AAABFFFFC0001440FFA9EACB005155401AE9C16B03AFE0;
defparam sp_inst_18.INIT_RAM_12 = 256'hE6C6C50FC0006FF905BA3A6A4DF54EA56A7774C6BC5BFFAFFBFABC000C000100;
defparam sp_inst_18.INIT_RAM_13 = 256'h2AC55AEAFFAFABFC003FC415003F1AA941F96954BE56AA5ABC03C000FC555038;
defparam sp_inst_18.INIT_RAM_14 = 256'h51A95AA955ABFFFF3FAC0555393FC6C4E5AF006FF9C5BCE4AAA1C3E955437729;
defparam sp_inst_18.INIT_RAM_15 = 256'h5AA5C17E4DAC6B3AA55394BB26E8555AABEABFFFFFC03FD55450FC6A941BE095;
defparam sp_inst_18.INIT_RAM_16 = 256'hFC3B013F154000C654C5BE45059155AA55555AFEABFFFFC054FE555B13D56F01;
defparam sp_inst_18.INIT_RAM_17 = 256'hAAABFCFFF0FAAFFFF000EBFBD546A9BF39F6CC4FFFAA600DA2EAC6956AAFAAFF;
defparam sp_inst_18.INIT_RAM_18 = 256'h3FAAA4D3DCEBCB6A96AAAAAFFFFFBD000C1A91546944BA55671AA55AA965555A;
defparam sp_inst_18.INIT_RAM_19 = 256'h0594563A55506AA5AAAA5555A5AAABFFFF3FBFEA555ABC153AFB06F8AB902BA3;
defparam sp_inst_18.INIT_RAM_1A = 256'hA550F1B5A93AAFD6936B3A20E3AA553A49881AFAAAAAAAAAFFFFFFC50F141530;
defparam sp_inst_18.INIT_RAM_1B = 256'h0FEAAAAABFFEAFFC153C53C3FF154147FA55546A96AAAA55555555AAFFFFFFFF;
defparam sp_inst_18.INIT_RAM_1C = 256'h656AAAA94040000556AAAAFAAA9553B215553C0F000E1C974EF9543940DC8FA3;
defparam sp_inst_18.INIT_RAM_1D = 256'h00F0392D3237903A4FE51D3AADC3FFFAABBFBEAC30000553B3055705456D6403;
defparam sp_inst_18.INIT_RAM_1E = 256'hFFC00F6503FDA411A54161A40546AAAA5550030FF0405556AAAAA94EC703F014;
defparam sp_inst_18.INIT_RAM_1F = 256'hFFC00000015555550FF7D56B03FFFF808958B0FF90E90E23AAB2BFAFEAAFFFFF;
defparam sp_inst_18.INIT_RAM_20 = 256'hA93940F9D25B15AAAFEAB0FFFFFFFC01540FCBE90B85364BA4651A6AA955500F;
defparam sp_inst_18.INIT_RAM_21 = 256'hF92900196E92A9A56AA565503FFC00033C000000143E95005AAAFEA4FE3EB16A;
defparam sp_inst_18.INIT_RAM_22 = 256'h3F03FF7BF11406A54FE40F11595E43C038DD6DA56AAFEAC0FCFFFBFF0515406F;
defparam sp_inst_18.INIT_RAM_23 = 256'h956AAA96C303FF0CFB0016459655A5051BAAABCF95AA555550FFFC15400FFFFF;
defparam sp_inst_18.INIT_RAM_24 = 256'hFBE5AA9505500FF05554003FFFFF03C6547043C030339FEC300394FC15274962;
defparam sp_inst_18.INIT_RAM_25 = 256'hFFFFB93929BE540FC167913E8AAAABAAAAFFC03C00F05015555016856A6ABFAB;
defparam sp_inst_18.INIT_RAM_26 = 256'h3003F1405150556E56BE96C2A9AC5AAAA5555503F1555400FBEBEBFC440C5FFF;
defparam sp_inst_18.INIT_RAM_27 = 256'h03C1555403EAAAAB14D044D5555A554E934153C0015549383F6AAAAAABEABF00;
defparam sp_inst_18.INIT_RAM_28 = 256'h1AAAA4D3E4F1BAAAAAAFAAB0C4FFFFC5500101A9BE96FEAB3A91A9AAAA9555A9;
defparam sp_inst_18.INIT_RAM_29 = 256'hA9BF47EBFA6AAA9AAEAA55AAA94015555503EAAFAC4F46E2AAAC03B2A40D0553;
defparam sp_inst_18.INIT_RAM_2A = 256'hABF0EA1BD9006FEAE5405ABEB9BC0E8E4F90C6AAAAAAAFFEBF10FABF000FF0A5;
defparam sp_inst_18.INIT_RAM_2B = 256'hAAAAAFFBFEF1403FFF00000555A5AA5A9AA58E9B1AFA5556AAAA555555540FAA;
defparam sp_inst_18.INIT_RAM_2C = 256'hA85AA9555AAAAA555555500FEAAF39A51F8E4063FFEA9A15A55300F92943E456;
defparam sp_inst_18.INIT_RAM_2D = 256'hC5690006FFFB910F93A5554A5A9AAABFFFFAC55400EB000550569696A56BEAEA;
defparam sp_inst_18.INIT_RAM_2E = 256'h5043EFFC1956AA6E55A5B0E55BA95AA5456AEAA55550100003EAFF815073F4D1;
defparam sp_inst_18.INIT_RAM_2F = 256'h55554000000FEBCD1541C54D24BC0EBEB0000F94E93FEAC0C9AA5AAAFFFF3F15;
defparam sp_inst_18.INIT_RAM_30 = 256'h53943C01C2FAAAAAAAFFFF01405001FFC06455BEF50AF47F9563F559A555ABE9;
defparam sp_inst_18.INIT_RAM_31 = 256'hBFD42F91AF2AEA9555A56AAAA9400500000003FF39A9076A93421A500014000E;
defparam sp_inst_18.INIT_RAM_32 = 256'hF0FFE42DBFE4E86A5A95500F39390FF0B1A6BEAAAAABFFFC143C0FF00FC191A6;
defparam sp_inst_18.INIT_RAM_33 = 256'hAABEAFFFF000F0FFB1400646957391FE9BB0FF1A5556956AAAA9400000000540;
defparam sp_inst_18.INIT_RAM_34 = 256'h72A55555A69A955000140415000003E5A2C0E4ED946A954FFBE4D3FC0B6CE07E;
defparam sp_inst_18.INIT_RAM_35 = 256'hC0EB69553A964E0F058700C63EFABEFFFEFC000FFFF51454C540B396FFAEFFF4;
defparam sp_inst_18.INIT_RAM_36 = 256'h43C3C556405600BEAFEF97EFE5A65500555A95555401696400400003E58BC0E7;
defparam sp_inst_18.INIT_RAM_37 = 256'h555405A95000010003EA1B00E0390B1410E8C4E401B1C553083FFAFFFFFAF0F1;
defparam sp_inst_18.INIT_RAM_38 = 256'h405CB1BF92A0FFEBFFFFEFC0C13F001955540406BFEABFEF9AAA05400015AAA5;
defparam sp_inst_18.INIT_RAM_39 = 256'h56FFA5BCFFABB9C00000556A95559555550000000000FC1BC3D4D3C6FFE9096E;
defparam sp_inst_18.INIT_RAM_3A = 256'h3000003016AFE4D55695038F5556DB6F039013FFAAFFFFFFCFF0F05555555054;
defparam sp_inst_18.INIT_RAM_3B = 256'hFFFABFEBFEFFC0C164065555A507BEA6FAF3FEAB00010555559596AA55540000;
defparam sp_inst_18.INIT_RAM_3C = 256'h9C0000400556AA9AAA95400000FF040000016FE503F93EA8AC15B2C6B0039FC3;
defparam sp_inst_18.INIT_RAM_3D = 256'hEA553E4FA3F06871AAF00F7540FFFAFFBFFAC01401502E40101562CBEBE6A83E;
defparam sp_inst_18.INIT_RAM_3E = 256'h03C030BA40405AFBEFEE5A6FA97FFAFFF0015696AAAA5000FC03F00400000C63;
defparam sp_inst_18.INIT_RAM_3F = 256'h55A5690000F05000500004FC6AA96950FE4FFFC72C3FC00E0643FFAFFEFFABC0;

SP sp_inst_19 (
    .DO({sp_inst_19_dout_w[29:0],sp_inst_19_dout[9:8]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[9:8]})
);

defparam sp_inst_19.READ_MODE = 1'b0;
defparam sp_inst_19.WRITE_MODE = 2'b00;
defparam sp_inst_19.BIT_WIDTH = 2;
defparam sp_inst_19.BLK_SEL = 3'b010;
defparam sp_inst_19.RESET_MODE = "SYNC";
defparam sp_inst_19.INIT_RAM_00 = 256'h3EAB869550155554395BFFAAAA55555555AAAA9A65AA9AAAEAAAAFAF00155555;
defparam sp_inst_19.INIT_RAM_01 = 256'hA9AAAAAAAAAAAAFEBC015555556AAAAA66AAAA556AA55550155A500015555554;
defparam sp_inst_19.INIT_RAM_02 = 256'hAAAAA9555555A9400C00000003EAAA1A550555543E6FFFFA55A955555556AAAA;
defparam sp_inst_19.INIT_RAM_03 = 256'h43FBC0F95555A9555555695AAAAAAAAAAAAAAAABFAB00155555AAAAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_04 = 256'hAFAAC055556AAAAAAAFAFAA5AAAAAAA5555556A903FBF00003FAAAADA9545555;
defparam sp_inst_19.INIT_RAM_05 = 256'hA40EAAFFCFFFEAAA86A55555540003FA955556A5555566956A9AAAAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_06 = 256'h5555556955AAAAAAAAAAAAAAAAAAAA056AAAFFFFFEAAAAAA55546AAAA555556A;
defparam sp_inst_19.INIT_RAM_07 = 256'hAAAAAAAAAAA9556AAAA55555AAA4EAAAFFFFFEBEA62AA555555540FE55555555;
defparam sp_inst_19.INIT_RAM_08 = 256'hE95DAA556555543EA555555555955555A55A9AAAAAAAAAAA6AAAAAA95555AAAA;
defparam sp_inst_19.INIT_RAM_09 = 256'hAAAAAAAAAAAAAAAAA5555555556AAAAAAAAAAAAAAAAAA95556AAA7EAAAAFFFAB;
defparam sp_inst_19.INIT_RAM_0A = 256'hAAAAAAAA555AAA93AAAAAAAAAA9586A55554143FA95555555555A555AA55A96A;
defparam sp_inst_19.INIT_RAM_0B = 256'hE9555555555556A55AA9AA55AAAAAAAAAAAAAAAAAA81555555555A9555555556;
defparam sp_inst_19.INIT_RAM_0C = 256'hAAAA155555555555A55555555555AAAAAA556ABE9E6AAAAAAAA9576A95550143;
defparam sp_inst_19.INIT_RAM_0D = 256'hFA4E56AAAAAA51B6AA5540140FA55555556A555AA5AAAAAA5AAAAAAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_0E = 256'h555AA9A9696AAAAAAAAAAAAAAAAAA9555555555556AA9555540005AAAAAAA5AA;
defparam sp_inst_19.INIT_RAM_0F = 256'h555AAAAA55550005AAAAAAAAAAAA4E55AA95A51B6AA5540543FA55555555AA55;
defparam sp_inst_19.INIT_RAM_10 = 256'hB5AA5555543E90015555556965556AA9A995AAAAAAAAAAAAAAAAAAA555555555;
defparam sp_inst_19.INIT_RAM_11 = 256'hAA9AAAAAAAAAAAAA95555555556AAAAAAA55550015AAAAAAAAAAAA5395A95555;
defparam sp_inst_19.INIT_RAM_12 = 256'h00156AA56AAAAAAA93959555571AA5555543EA5001555555555556AAA6AAAAAA;
defparam sp_inst_19.INIT_RAM_13 = 256'h4015555555555556AA956AAAAA95AAAAAAAAAAAAAA55555556A96AAA56AAAA95;
defparam sp_inst_19.INIT_RAM_14 = 256'hAAA95555555555559556AAAA9540156A5555AAAAAA5396555561695555543E95;
defparam sp_inst_19.INIT_RAM_15 = 256'hAAAA53955156C595555400E94001555555555555556A956AAAAA56AAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_16 = 256'h5695AA95AAAAAA6AAA6AAAAAAAAAA555555555555555556AAA555555A95555AA;
defparam sp_inst_19.INIT_RAM_17 = 256'h555556555A5555555AAA55556AAAAA4E950568655555400FA900155555555555;
defparam sp_inst_19.INIT_RAM_18 = 256'h95555503FA55505555555555555556AAA6AAAAAAAAAAAAAAA9AAAA9555555555;
defparam sp_inst_19.INIT_RAM_19 = 256'hAAAAAAEAAAAAAAAA555555555555555555955555555556AA9555AAAA4E5555B5;
defparam sp_inst_19.INIT_RAM_1A = 256'h5555055AAA95556AA94E95AC195555400FA55555555555555555556AA5AAAA9A;
defparam sp_inst_19.INIT_RAM_1B = 256'hA555555555555556AA96A96955AAAAAAAAAAAAAAA95555555555555555555555;
defparam sp_inst_19.INIT_RAM_1C = 256'hAAA55555555555555555555555555405AAAA96A5AAA54FAAC155554000FA5005;
defparam sp_inst_19.INIT_RAM_1D = 256'hAA5A954FEF0555400FFFE54001695555555555569AAAAAA959AAA9AAAAAAAAA9;
defparam sp_inst_19.INIT_RAM_1E = 256'h556AA5AAA956AAAAAAAAAAAAAAAA955555555450055555555555555015A95AAA;
defparam sp_inst_19.INIT_RAM_1F = 256'h001555555555555550055555A95555550FFC050000FFFA940005555555555555;
defparam sp_inst_19.INIT_RAM_20 = 256'h003FFFAA5400555555555A55555556AAAAA56AAAAAAA9AAAAAAAAA5555555550;
defparam sp_inst_19.INIT_RAM_21 = 256'hAAAAAAAAAAAAAAA95555555540015554415555555540155555555555003FF000;
defparam sp_inst_19.INIT_RAM_22 = 256'h405400400555555550000F00000FFEBFEA5001555555556A56555555AAAAAAAA;
defparam sp_inst_19.INIT_RAM_23 = 256'h5555555569A955A655AAAAAAAAAAAAAAAAAAAABAA55555555500015555500000;
defparam sp_inst_19.INIT_RAM_24 = 256'hAA9555555555500555555540000054140005541545440FFC3003FFABFFE95005;
defparam sp_inst_19.INIT_RAM_25 = 256'h0000003FFFFFFFFABFFEA9401555555555556A96AA5AAAAAAAAAAAAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_26 = 256'h9AA95AAAAAAAAAAAAAAAAABEAAAB5555555555540555555500000001500C0000;
defparam sp_inst_19.INIT_RAM_27 = 256'h5415555554000000550000C00000000FFEFFFEBFFFFFFA9540555555555555AA;
defparam sp_inst_19.INIT_RAM_28 = 256'hFFFFFFA9550555555555555A6A55556AAAAAAAAAAAAAAAAAEAAAA95555555555;
defparam sp_inst_19.INIT_RAM_29 = 256'hAAAAAAAAAAAAAAA555555555555555555554000001500003FFFC03F3FFFBFFFE;
defparam sp_inst_19.INIT_RAM_2A = 256'h000500000FFFFFFFFFFFFFFFFFFC0FFAA55515555555555555AA5555AAA55AAA;
defparam sp_inst_19.INIT_RAM_2B = 256'h55555555555AAA9555AAAAAAAAAAAAAAAAAABAAAD55555555555555555555000;
defparam sp_inst_19.INIT_RAM_2C = 256'hAB555555555555555555555000004000000FFFF3FFFFFF00000300FFEAA95555;
defparam sp_inst_19.INIT_RAM_2D = 256'hC00000000000000FFEAAAAA55555555555556AAAAA55AAAAAAAAAAAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_2E = 256'hAAA95556AAAAAAAAAAAAAFAAAAA95555555555555555555554000000000400FF;
defparam sp_inst_19.INIT_RAM_2F = 256'h5555555555500010000015503C01500005555000FFEAAABFA5555555555595AA;
defparam sp_inst_19.INIT_RAM_30 = 256'h03FFEBFFC3955555555555AAAAAAAA556AAAAAAAAAAAAAAAAAAEA55555555555;
defparam sp_inst_19.INIT_RAM_31 = 256'hAAAAAAAAAAEAAA95555555555555555555555400400000555400555555555550;
defparam sp_inst_19.INIT_RAM_32 = 256'h050000015555015555555550403FFAAFF003955555555556AA96A55AA56AAAAA;
defparam sp_inst_19.INIT_RAM_33 = 256'h555555555AAA5A555AAAAAAAAAAEAAAAAAAFAAAA555555555555555555555555;
defparam sp_inst_19.INIT_RAM_34 = 256'hAD555555555555555555555555555400056A5501555555500000FEABFF010395;
defparam sp_inst_19.INIT_RAM_35 = 256'h1500555540000FFAFFC0550E955555555556AAA5555AAAAA6AAAAEAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_36 = 256'hA9696AAAAAAAAAAAAAAAAAAAAAA5555555555555555555555555555400156A54;
defparam sp_inst_19.INIT_RAM_37 = 256'h5555555555555555540055AA554000555500C0FFFFF015543A95555555555A5A;
defparam sp_inst_19.INIT_RAM_38 = 256'hFFFC055554EA55555555556A6A95AAAAAAAAAAAAAAAAAAAAAAAA955555555555;
defparam sp_inst_19.INIT_RAM_39 = 256'hAAAAAAABAAAAAA1555555555555555555555555555550155695503C000000FFF;
defparam sp_inst_19.INIT_RAM_3A = 256'h4555554555555500000003FAFFFFC055A954E95555555555655A5AAAAAAAAAAA;
defparam sp_inst_19.INIT_RAM_3B = 256'h5555555555556A6AAAAAAAAAAAAAAAAAAAAEAAA8555555555555555555555555;
defparam sp_inst_19.INIT_RAM_3C = 256'hA15555555555555555555555550055555555555554003FFFABFFF0155AA953A9;
defparam sp_inst_19.INIT_RAM_3D = 256'h5555400FFEAFFC05555AA543AA55555555556AAAAAAAAAAAAAAAAEBAAAAAABEA;
defparam sp_inst_19.INIT_RAM_3E = 256'hA96A9AAAAAAAAAAAAAAAAAAAAA80000005555555555555550154055555555159;
defparam sp_inst_19.INIT_RAM_3F = 256'h55555555550555555555550155555555000FFFC056956AA54EA955555555556A;

SP sp_inst_20 (
    .DO({sp_inst_20_dout_w[29:0],sp_inst_20_dout[11:10]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[11:10]})
);

defparam sp_inst_20.READ_MODE = 1'b0;
defparam sp_inst_20.WRITE_MODE = 2'b00;
defparam sp_inst_20.BIT_WIDTH = 2;
defparam sp_inst_20.BLK_SEL = 3'b010;
defparam sp_inst_20.RESET_MODE = "SYNC";
defparam sp_inst_20.INIT_RAM_00 = 256'h48AA377F755DFDF76000808828A0AA8A80080000000A82A2028200A0DDF5FFFD;
defparam sp_inst_20.INIT_RAM_01 = 256'h00008202800228028177557D7FD5FFF5FFD5FFD7D57D5FD5FFDDF57D755FFFFD;
defparam sp_inst_20.INIT_RAM_02 = 256'hDD7FDD75D5FDFDFDD1F557FD74802875F75F7FDF4802A0A282200A082AA000A8;
defparam sp_inst_20.INIT_RAM_03 = 256'hDE08158A882080A0AAAA828220A2082A82AA80080087DF55FD555575FD7FD77D;
defparam sp_inst_20.INIT_RAM_04 = 256'h000AB5F57F57F555555757D5FF5F5F75D5F7F7FDDC2225D7D480A0A15FD5D5FD;
defparam sp_inst_20.INIT_RAM_05 = 256'h5550022812288022B55FFD57DF7D5EA08000A80AAA8A000A2A822AAAAAA2AA08;
defparam sp_inst_20.INIT_RAM_06 = 256'h0AAA2A00A82828282AA00A82A0A8A85DD5F57FFFF57D7DFD755D57F7D7D5D7DF;
defparam sp_inst_20.INIT_RAM_07 = 256'hD5FFFF5F7FDDD7DDF7F5D5FDD577200280A02AA80AFD5F5FDD5F7D888820A2AA;
defparam sp_inst_20.INIT_RAM_08 = 256'h800177FFFDD57FC0A0220AAAAA0AAA888A8082A8A0AA8A8A08808281557F57FF;
defparam sp_inst_20.INIT_RAM_09 = 256'hAA008AA202800820055FF555FF55555F757FDFD77DFF5DFFF77D5E8028A80A8A;
defparam sp_inst_20.INIT_RAM_0A = 256'h55F557575FDDFFF400A00AA0082A17F5D7D777E8A20020AAAAA802AA2A28008A;
defparam sp_inst_20.INIT_RAM_0B = 256'hA88AA280AAAAA80282000828222AA00A8088202A2A17FD5555FFD557FFD55557;
defparam sp_inst_20.INIT_RAM_0C = 256'h0AAA7D7FD5FFFFF557FFD57FD7D5D555575F77FD7A8880002A2800F5D55DDFFC;
defparam sp_inst_20.INIT_RAM_0D = 256'hFFF80A80200022877F57777D5A2802A800082AA0080A8008A20AAA802080A8A0;
defparam sp_inst_20.INIT_RAM_0E = 256'hA020000022A0A228A8020082A000295FF5FFF55FD57D75F57D7FFD55F5D5F5F7;
defparam sp_inst_20.INIT_RAM_0F = 256'h5557FF55FD7D757F57F55D7FF7F77020A822A008D5D5775FD42A208A8000A88A;
defparam sp_inst_20.INIT_RAM_10 = 256'h8DD75F5F75682AA80200AA2002AA800020082A2AA220A828028280A5FFD55555;
defparam sp_inst_20.INIT_RAM_11 = 256'hAA0AA80A8000AAAA17FFFD55557D57FDD55F5777DFFF5D557FFD57DE0A0202AA;
defparam sp_inst_20.INIT_RAM_12 = 256'hDDDDF5F57FFFD7F776A8A282A0DDDFF55D542200AA080AA8082AA8A000002A00;
defparam sp_inst_20.INIT_RAM_13 = 256'hA2800AAA02AAAAA000000AAA2A00200080A2A08A2A5FFFFFD55555555DFFF575;
defparam sp_inst_20.INIT_RAM_14 = 256'h2A015FFD57FD555D57FD5FFF777FF7777FF5F5D55DF6A220AA8F7DF5557742AA;
defparam sp_inst_20.INIT_RAM_15 = 256'hFF7DDE28AAAAB55FF55DD7802828000AA82A2AAAAA800AAAAAA822802AA28208;
defparam sp_inst_20.INIT_RAM_16 = 256'h002AAA0A20A0AA002A0A28AA080AA5FF55555FFFFF5FFF55F5FDF55DDF757D57;
defparam sp_inst_20.INIT_RAM_17 = 256'hFFFD557F55FD55555FFF7D7F7F57DD5888A82BF57FFFFFF2AA0A82802AAAAA08;
defparam sp_inst_20.INIT_RAM_18 = 256'hFDF7F5DC8A28A82A02AAAAA8A20AA28000A02AA882AA280A88200297F575577F;
defparam sp_inst_20.INIT_RAM_19 = 256'hAA0AA828AA2A8000FFFF5555FFFFFFFFFD5FFFF7FFFF55FF7FFF575D7202A005;
defparam sp_inst_20.INIT_RAM_1A = 256'h5FF5FDDD575D7FDFF7F28283FDFD55DF78AA8AA8AAAA28AA8AAAAA0A882A2082;
defparam sp_inst_20.INIT_RAM_1B = 256'h082AAA22A82AAA00AA22080080AA8AA2A8AAA88003FFFD5555555557FFFFFFFF;
defparam sp_inst_20.INIT_RAM_1C = 256'h8A0FFFF5557FFFF555555FFFFD5FF75FFF7F555F5D7D588ABF5D57DD7F02880A;
defparam sp_inst_20.INIT_RAM_1D = 256'h57FFFF7A22FDDFDF7820008022A8000A8AA2AA2000282AA2802AA82AA80A8A80;
defparam sp_inst_20.INIT_RAM_1E = 256'hA0002082008208220A8A0A0A28809FFF5557FFFF7FFFFFF5555557DD755555FD;
defparam sp_inst_20.INIT_RAM_1F = 256'hF7FFFDFDFFD57FFFDFF7D55D55FFFD55F229775DD70A22A0A82200202AA2A0AA;
defparam sp_inst_20.INIT_RAM_20 = 256'hD5C20A882AA8A0AAA02A80082AAA00022A200282802A0802088A8A57FD5557FF;
defparam sp_inst_20.INIT_RAM_21 = 256'h02000A2AA808020157555557FFFFFFF55577FFF57D5D57FF55D5FD5DFDC28F57;
defparam sp_inst_20.INIT_RAM_22 = 256'h5555775D5DFF5D5FDFDFD0FFFD5882AA880222202AA02A2A20AAAA80AA2A828A;
defparam sp_inst_20.INIT_RAM_23 = 256'h202AAA82002828002A28A08A28AA0AA2A20000AA2555555557FFFFF5FFD55555;
defparam sp_inst_20.INIT_RAM_24 = 256'hA2155755D557FFFF575FF555555D55D7575FFD55757770A1455620AA80802028;
defparam sp_inst_20.INIT_RAM_25 = 256'hFFF77D4828A8AA0A8020AAAA8AAAA8AAAA800A228882A0A2AAA8A82A80800A02;
defparam sp_inst_20.INIT_RAM_26 = 256'h00000AA2AA22AA8028202888000855575555557F7FF57FFF557FFF557551F555;
defparam sp_inst_20.INIT_RAM_27 = 256'h7FFF555FFD55FFFF55755795555F57F2A208080000A88A28A082AAAAA82A800A;
defparam sp_inst_20.INIT_RAM_28 = 256'h200028220A0202AAAAA0AA800A20808AAA0AAA222A28A000200A01555555557D;
defparam sp_inst_20.INIT_RAM_29 = 256'h022A2A82A08800057D555555F55FD5557FF57FFFFDDDD77E0A83FC0C200800A8;
defparam sp_inst_20.INIT_RAM_2A = 256'hFFF5F5575200220808000A8AA22BF0888A220A2AAAAAA28280A8AAA82A00820A;
defparam sp_inst_20.INIT_RAM_2B = 256'hA2AAA00A0A82A80A0820002AAA0A00000208882217FD555557F55555555FD57F;
defparam sp_inst_20.INIT_RAM_2C = 256'h0A57F55F57FFFD555557FF557FFD75577FD8800E0A0AA85F5DDE7F888A822008;
defparam sp_inst_20.INIT_RAM_2D = 256'h15FDFFFDFFD57570A20AAA022A82AA80200A0AAA002A002AAA0020200A8A8080;
defparam sp_inst_20.INIT_RAM_2E = 256'h2AA02A0022A000A8A00A208AA2035555FD5FFFF555575FFFF57F757F7D5F5F20;
defparam sp_inst_20.INIT_RAM_2F = 256'h55557FFFFFF57D5DFFD555F7EB77D7FFF555FDD5820A828202AA0AAA800A08AA;
defparam sp_inst_20.INIT_RAM_30 = 256'hDCA8200A3EAAAAAAAA82080A82A00228088AAA28A2A0A2AA2A822F5555D55FFF;
defparam sp_inst_20.INIT_RAM_31 = 256'hA8A8AA020A02803FFD55555FFD5FF5FFFFFFF55555555D7D7D7F757FF57D55F5;
defparam sp_inst_20.INIT_RAM_32 = 256'h557FF55D5F777D75757FF5FFF762000227FC82AAAAAA2828AA00080002020208;
defparam sp_inst_20.INIT_RAM_33 = 256'hAAA2A808A2A02022828028882A202AA82220AAA0D7F5555557FD5FFFFFFFFFFD;
defparam sp_inst_20.INIT_RAM_34 = 256'hA955F7FD5557D55FFFFFFFFFFD5555DF55FF7F755FD57FDFD5772020A2D7F602;
defparam sp_inst_20.INIT_RAM_35 = 256'h5F7DD7FF757DD880289FDF7A820A82A00A808000020AAAA82A820222AA00AAA2;
defparam sp_inst_20.INIT_RAM_36 = 256'hA0028AA8A2AA822A2A082AAA80057FFFF555555557FF5557FFFFD557DF7FFF75;
defparam sp_inst_20.INIT_RAM_37 = 256'h5555FDF55FFFFFD555F5F5DF7FDD57FD7755958A28ADDFFDCA800A02802A0202;
defparam sp_inst_20.INIT_RAM_38 = 256'hAA8B77557D2A00280200AA080A80A822A2AA2808A8002A8A00001FFFDFFD5FD5;
defparam sp_inst_20.INIT_RAM_39 = 256'hA0A00028AA00285F5FFFFD5F5555555555FFFFFFD555FF7DFF77DC375FF75228;
defparam sp_inst_20.INIT_RAM_3A = 256'h5557D5757F5577D5557F560082823DDFFF7F0800AAA80200000802AAAAAAA088;
defparam sp_inst_20.INIT_RAM_3B = 256'h02AAA0280A800A0A8808AAAA0AAA2A80A8A02829555FFFFD555557FD5F5FDFFF;
defparam sp_inst_20.INIT_RAM_3C = 256'h0D555FFFFF55F55FFF5FFF55FD557FF55555F775F57F4800A2808DFF7D5F5480;
defparam sp_inst_20.INIT_RAM_3D = 256'h7F55DF72802A297555FFFD5EA8002A82A02A0A820AA00880AAAA888A22808028;
defparam sp_inst_20.INIT_RAM_3E = 256'hA002022080A2A0A0882A000A02BFFF5557FF55D5FD7F7FFF57FD557FD5557DDD;
defparam sp_inst_20.INIT_RAM_3F = 256'h55555DFFFD57FFFFFD5555FDD7FD7D7F5F50A837DDFFFFFFFAA802A02A80A82A;

SP sp_inst_21 (
    .DO({sp_inst_21_dout_w[29:0],sp_inst_21_dout[13:12]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[13:12]})
);

defparam sp_inst_21.READ_MODE = 1'b0;
defparam sp_inst_21.WRITE_MODE = 2'b00;
defparam sp_inst_21.BIT_WIDTH = 2;
defparam sp_inst_21.BLK_SEL = 3'b010;
defparam sp_inst_21.RESET_MODE = "SYNC";
defparam sp_inst_21.INIT_RAM_00 = 256'h4FAA8F3FEAABFA54D3AD690FEA5A55656AAAAAAAAAAAAAAF3FFEF0F06BF00001;
defparam sp_inst_21.INIT_RAM_01 = 256'hAAAAAAAABFFFEB03C2AF000140155555001500FF15400FFABFC0EA96AFFAAAAA;
defparam sp_inst_21.INIT_RAM_02 = 256'h01555030FFFC0096555AAAAA94FA9670FEAAFFA434C55A5255AAA556955AAAAA;
defparam sp_inst_21.INIT_RAM_03 = 256'h5E91BF9E515AAA555555696AEAAAAAAAAAAABFFC0FCABF000155555A55555455;
defparam sp_inst_21.INIT_RAM_04 = 256'hF0FFEFF000555AAAAAA9A9500055A540C0F3F003553F0569650FAA5E0FFABFFA;
defparam sp_inst_21.INIT_RAM_05 = 256'h5253FF015440FFE94C0FEBFEA43C0E43A55556A55565AAA5AAAAEAAAAAAAAAAB;
defparam sp_inst_21.INIT_RAM_06 = 256'hA55595AA56AAABEBEAAFFAAAAFFFFFFC155AAAAAAA9541553FFAC55953FFC3C0;
defparam sp_inst_21.INIT_RAM_07 = 256'h6A5555559550FFC15940FFFC154D3FFFC0003FFF91700FFFFAA54FA3A5455555;
defparam sp_inst_21.INIT_RAM_08 = 256'hF90A03FFFFAA94E4EA94555555A55566A56AAAABAFAABFFAABBFFFFC00005555;
defparam sp_inst_21.INIT_RAM_09 = 256'hAAFFAAAFFEBFFBEFF00FF0000055555555555014015550FFF05548FFFFFC0FFF;
defparam sp_inst_21.INIT_RAM_0A = 256'h550555540FC15538FFFFFFFFFF8F4C3FFFF954E53EAA95555556A955AA96AA6A;
defparam sp_inst_21.INIT_RAM_0B = 256'h4FA5556A555556A96AFAAA96AAEAAFFABFBFEFEAAAFFFC000000155400000000;
defparam sp_inst_21.INIT_RAM_0C = 256'hFAAAFC00000000055400003FFFC01555540F0555226BFFFFEAE4F3B0FFFA554F;
defparam sp_inst_21.INIT_RAM_0D = 256'h54DE56BFEAAA7F3B3FFE9455393AA956AAAA955AA6AAAAAA5AEAAABFEFBFFFAF;
defparam sp_inst_21.INIT_RAM_0E = 256'h5A9AAAAAA96FAAEAABFEFFFEAFFFE80005000550155545003FEAAC5505550005;
defparam sp_inst_21.INIT_RAM_0F = 256'h55555555003FEAAC540555400554D246AB9554F370FFE9555393EAA56AAAAA65;
defparam sp_inst_21.INIT_RAM_10 = 256'h37C3FAA5A925240155AA55AAA9556AAAAAA6AAAAAAAFFBEBFEBEBFA000155555;
defparam sp_inst_21.INIT_RAM_11 = 256'hAAAAABFABFFFAABFC000015555555555555003EABC005155400154E391A9554F;
defparam sp_inst_21.INIT_RAM_12 = 256'hA6BC05000000155427915414377CFAAAAA9383E00056A556A69556AAAAAAAAAA;
defparam sp_inst_21.INIT_RAM_13 = 256'h40155555A955555AAAAAAAAAAAAAAFFFABFEBFBAFF0000001555555551555543;
defparam sp_inst_21.INIT_RAM_14 = 256'hEAFC0000000155515401555543EAAF043FF0001550E795400022FFAAAA9438EA;
defparam sp_inst_21.INIT_RAM_15 = 256'h0040E3953C01DFFAAAA503938141555556955555556AA56AAAAA9ABFEAAFFAFB;
defparam sp_inst_21.INIT_RAM_16 = 256'hAA95AAA5AFAAAAAFEAAAFFAAABFAA00000000000005000555500FFFC103FFC00;
defparam sp_inst_21.INIT_RAM_17 = 256'h000155405500000000003C3F000010E350F158BFEAAA4FFD0E501555555555A6;
defparam sp_inst_21.INIT_RAM_18 = 256'hEBAAA90FA3EB91555555555659A55AAAAAAFEAAABEAAFFFABAAFFE8000000000;
defparam sp_inst_21.INIT_RAM_19 = 256'hAAFAAB3FAAEABFFF000000000000000001500003FFFF00003FFF0050D243C58B;
defparam sp_inst_21.INIT_RAM_1A = 256'h0FFFABC1540FFFC00392546C6FAAAA503A396AAA55555555655555AAA6AAAFAA;
defparam sp_inst_21.INIT_RAM_1B = 256'hFA955555569555AAAA9AFAAA6AAAAAAFFFAAAABFFC0000000000000000000000;
defparam sp_inst_21.INIT_RAM_1C = 256'hBAF00000003FFFF000000000000FFEAB0040000F0C3F93A6C6FAA9503FE7A556;
defparam sp_inst_21.INIT_RAM_1D = 256'h03FFFA93EF1BA5503FEA4E5545AAAAA55559555AAAAAAAA96AAAAAAAABFEBAAA;
defparam sp_inst_21.INIT_RAM_1E = 256'h5AAAAABEAA6AFAAAFAAAFAFAABAFC0000003FFFFFFFFFFF0000003FAAC000000;
defparam sp_inst_21.INIT_RAM_1F = 256'hFFFFFFFFFFC03FFFFAAFFFFC00FFFFEA43FC595503FA94E90145AA9A95595A55;
defparam sp_inst_21.INIT_RAM_20 = 256'h14FEA550E40155555A956AA69555AAAAEAAAAFFEAFEAABEFFABABF00000003FF;
defparam sp_inst_21.INIT_RAM_21 = 256'hFEBFAAAABFFBFEFC00000003FFFFFFFFFFFFFFFFFFFABEAAFFFFFFFA5503C054;
defparam sp_inst_21.INIT_RAM_22 = 256'hFFFFEAE6ABAAABFAA5500000000FA95550E40595555A95AA9A55556AAAAAAABF;
defparam sp_inst_21.INIT_RAM_23 = 256'h95555555AAAA96AA95AAAFAAEBAAFAAEAFFFFFFFE000000003FFFFF0FFFFFFFF;
defparam sp_inst_21.INIT_RAM_24 = 256'hFF000000C003FFFF030FFFFFFFFBFFBD546AAAAA9A9940F00003EA556A539406;
defparam sp_inst_21.INIT_RAM_25 = 256'h5559550FFFFFAAA56AA90E5415555655556AAA9AAA6AAAAEAAAAABEABFBFFFFF;
defparam sp_inst_21.INIT_RAM_26 = 256'hAAAAAAAAAAEAAABFEBFFEBCFFFFC00000000003FFFF03FFFFFEAAAFFE5515AAA;
defparam sp_inst_21.INIT_RAM_27 = 256'h3FFF000FFFFFAAAAFF95541555555403FEFBFAAAAAAAA03A5569555556956AAA;
defparam sp_inst_21.INIT_RAM_28 = 256'hAFFFEA43F955A955555A556AAA9A6A6AAAAAAAFEFFEBFFFF3FFAFC0000000000;
defparam sp_inst_21.INIT_RAM_29 = 256'hFEFFEBFFFFBFFFF000000000000FC0003FFFEAAAABFA55930FC000003FFBFFAA;
defparam sp_inst_21.INIT_RAM_2A = 256'hAAAFAA5A93FFF00C0FFFFFCFFEFFFFA50FE95595555559696AAA5556AAAA6AFA;
defparam sp_inst_21.INIT_RAM_2B = 256'h55555AA5A56AAAA5A6AAAAAAAAFAFFFFFFFBCFEF0000000000000000000FFFEA;
defparam sp_inst_21.INIT_RAM_2C = 256'hFF00000F000000000003FFFFEAABEAA95A50FFC0000FFC10500F3FFA5003E956;
defparam sp_inst_21.INIT_RAM_2D = 256'h155500015555403FA95000395555556A9AA5AAAAAA95AAAAAAFFEFEFFABFFFFF;
defparam sp_inst_21.INIT_RAM_2E = 256'hEAAA95AAAEAFFFBFAFFAF0FAAFFF0000FC00000000030FFFFFEAEF95956AA43F;
defparam sp_inst_21.INIT_RAM_2F = 256'h00003FFFFFFFEBFA5555BFE93C5AA9555AAA5500FEA55569795555556AA5A6AA;
defparam sp_inst_21.INIT_RAM_30 = 256'h0FAA9AAAFE2555555569A6AAAAAAAA96AABAAAFFFEAFFEBFEAB3FF0000C00000;
defparam sp_inst_21.INIT_RAM_31 = 256'hFCEABFFAFF3FFFFFFC000000000FF0FFFFFFFFFFFAAA56FC3A41AFEAAAAAAA55;
defparam sp_inst_21.INIT_RAM_32 = 256'hFFEAA96B003E96FFEFEAAA55543EAAAAF00EE95555559696AAAAA6AAA9AAFAFB;
defparam sp_inst_21.INIT_RAM_33 = 256'h555956A65AAA9A996AAAABABEAF0EAFFEFF0FFAFC3F0000000000FFFFFFFFFFF;
defparam sp_inst_21.INIT_RAM_34 = 256'hBC00F3FC0000000FFFFFFFFFFFFFFFA5AC003E9BFABFEAA55543EA9AAF154CE9;
defparam sp_inst_21.INIT_RAM_35 = 256'hAA96BEAA95410FAAABC16577A9A5695AA56AAAAAA9AAAAAAAAAAC3EFFFFFFFFE;
defparam sp_inst_21.INIT_RAM_36 = 256'hAAA96AABAAAAAAFFFFFFEBFFFFF03FFFF000000003FF0003FFFFFFFEA5AC003E;
defparam sp_inst_21.INIT_RAM_37 = 256'h0000FC000FFFFFFFFFAAB0103AA505AAA954C0FAABF16AA5DEAAA5A96A95AAAA;
defparam sp_inst_21.INIT_RAM_38 = 256'hAABC5AFFE4BAAA96A9AA55AAAAAAAAAEAEAAAAABFC3FFFFFFFFFBFFFFFFC0000;
defparam sp_inst_21.INIT_RAM_39 = 256'hAFF0FFFCFFFFFFFFFFFFFC000000000000FFFFFFFFFFAAFC003E5005A5540EFF;
defparam sp_inst_21.INIT_RAM_3A = 256'hFFFFFFEFFF003E55554003EABEBF06BFFFE77AAA5556A9AAAAAAAAAAAAAAAABA;
defparam sp_inst_21.INIT_RAM_3B = 256'hA9555A96A56AAAAABAABAAAAFAABFFFFFFF03FFFFFFFFFFC000000000F0FFFFF;
defparam sp_inst_21.INIT_RAM_3C = 256'hFBFFFFFFFF000000000FFFFFFFFFFFFFFFFFF03FAA940FFE5ABFC16AFC0FE73A;
defparam sp_inst_21.INIT_RAM_3D = 256'h3FFFA543FAAAFC5BFFFFFF9DEAAA95695A95AABEAAAABFAAAAAABFCF3FFFFC3F;
defparam sp_inst_21.INIT_RAM_3E = 256'hAAAAAAFFAAAAAFFFFC3FFFFFFEAAAAFFFFFF000000003FFFFFFFFFFFFFFFEBC0;
defparam sp_inst_21.INIT_RAM_3F = 256'h000000FFFFFFFFFFFFFFFFABC3FFFFEAA540FC05BCFFFFFE77AAA95A956A56AA;

SP sp_inst_22 (
    .DO({sp_inst_22_dout_w[29:0],sp_inst_22_dout[15:14]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,ad[14],ad[13]}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:14]})
);

defparam sp_inst_22.READ_MODE = 1'b0;
defparam sp_inst_22.WRITE_MODE = 2'b00;
defparam sp_inst_22.BIT_WIDTH = 2;
defparam sp_inst_22.BLK_SEL = 3'b010;
defparam sp_inst_22.RESET_MODE = "SYNC";
defparam sp_inst_22.INIT_RAM_00 = 256'hA5556AEAAAAAAAAA5401555000000000000000000000000040000505AAAFFFFF;
defparam sp_inst_22.INIT_RAM_01 = 256'h000000000000005416AAFFFFFFFFFFFFFFFFFFAAFFFFFAAAAABFAAAAAAAAAAAA;
defparam sp_inst_22.INIT_RAM_02 = 256'hFFFFFFEFAAABFFAAAAAAAAAAAA5555AFAAAAAAAA951555540000000000000000;
defparam sp_inst_22.INIT_RAM_03 = 256'hA555555000000000000000000000000000000001501AAAFFFFFFFFFFFFFFFFFF;
defparam sp_inst_22.INIT_RAM_04 = 256'h05002AAFFFFFFFFFFFFFFFFFFFFFFFFFBFAEAFFEAA95AAAAAAA55556FAAAAAAA;
defparam sp_inst_22.INIT_RAM_05 = 256'hFEA955AAAAAA55556BFAAAAAAA96A55400000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_06 = 256'h000000000000000000000000000000ABFFFFFFFFFFFFFFFFEAAABFFFFEAABEBF;
defparam sp_inst_22.INIT_RAM_07 = 256'hFFFFFFFFFFFFAABFFFFFAAABFFFA95556AAA955555AFFAAAAAAAA55400000000;
defparam sp_inst_22.INIT_RAM_08 = 256'h5556FEAAAAAAAA550000000000000000000000000000000000000003FFFFFFFF;
defparam sp_inst_22.INIT_RAM_09 = 256'h00000000000000000FFAAFFFFFFFFFFFFFFFFFFFFFFFFFAAAFFFFA555556A555;
defparam sp_inst_22.INIT_RAM_0A = 256'hFFFFFFFFFABFFFEA5555555555506BEAAAAAAA55400000000000000000000000;
defparam sp_inst_22.INIT_RAM_0B = 256'h5000000000000000000000000000000000000000002AABFFFFFFFFFFFFFFFFFF;
defparam sp_inst_22.INIT_RAM_0C = 256'h0000ABFFFFFFFFFFFFFFFFEAAABFFFFFFFFAFFFFE9555555555505AFAAAAAAA5;
defparam sp_inst_22.INIT_RAM_0D = 256'hFFA555555555405AEAAAAAAA9540000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_0E = 256'h000000000000000000000000000003FFFFFFFFFFFFFFFFFFEAAAABFFFFFFFFFF;
defparam sp_inst_22.INIT_RAM_0F = 256'hFFFFFFFFFFEAAAABFFFFFFFFFFFFA95555555505AFAAAAAAA954000000000000;
defparam sp_inst_22.INIT_RAM_10 = 256'h5ABEAAAAAA954000000000000000000000000000000000000000000FFFFFFFFF;
defparam sp_inst_22.INIT_RAM_11 = 256'h00000000000000003FFFFFFFFFFFFFFFFFFFFEAAABFFFFFFFFFFFFA955555550;
defparam sp_inst_22.INIT_RAM_12 = 256'hAAABFFFFFFFFFFFFE955555545ABAAAAAAA95400000000000000000000000000;
defparam sp_inst_22.INIT_RAM_13 = 256'h000000000000000000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFE;
defparam sp_inst_22.INIT_RAM_14 = 256'h0003FFFFFFFFFFFFFFFFFFFFFEAAAAFFEAAFFFFFFFA95555555AAAAAAAAA9500;
defparam sp_inst_22.INIT_RAM_15 = 256'hFFFFA95541556AAAAAAAA9540000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_16 = 256'h00000000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFAAABFFEAABFF;
defparam sp_inst_22.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFEBEAFFFFFFA9550556AAAAAAA5555000000000000000;
defparam sp_inst_22.INIT_RAM_18 = 256'hAAAAAAA554000000000000000000000000000000000000000000003FFFFFFFFF;
defparam sp_inst_22.INIT_RAM_19 = 256'h0000004000000000FFFFFFFFFFFFFFFFFFFFFFFEAAAAFFFFEAAAFFFFA954156A;
defparam sp_inst_22.INIT_RAM_1A = 256'hFAAAAABFFFFAAABFFEA95556AAAAAAAA95400000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1B = 256'h000000000000000000000000000000000000000003FFFFFFFFFFFFFFFFFFFFFF;
defparam sp_inst_22.INIT_RAM_1C = 256'h000FFFFFFFEAAAAFFFFFFFFFFFFAAAAAFFFFFFFAFBEAA9556AAAAAAA95540000;
defparam sp_inst_22.INIT_RAM_1D = 256'hFEAAAAA955AAAAAA955550000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_1E = 256'h00000000000000000000000000003FFFFFFEAAAAAAAAAAAFFFFFFEAAABFFFFFF;
defparam sp_inst_22.INIT_RAM_1F = 256'hAAAAAAAAAABFEAAAAAAAAAABFFAAAAAAA956AAAAA95555000000000000000000;
defparam sp_inst_22.INIT_RAM_20 = 256'hAA5555550000000000000000000000000000000000000000000000FFFFFFFEAA;
defparam sp_inst_22.INIT_RAM_21 = 256'h0000000000000003FFFFFFFEAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA96AAA;
defparam sp_inst_22.INIT_RAM_22 = 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAA5555555000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_23 = 256'h00000000000000000000000000000000000000000FFFFFFFFEAAAAAFAAAAAAAA;
defparam sp_inst_22.INIT_RAM_24 = 256'h007FFFFFBFFEAAAAFEFAAAAAAAAAAAAAAAAAAAAAAAAAAA5AAAA9555555540000;
defparam sp_inst_22.INIT_RAM_25 = 256'hAAAAAAA555555555555550000000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_26 = 256'h0000000000000000000000100001FFFFFFFFFFEAAAAFEAAAAAAAAAAAAAAAAAAA;
defparam sp_inst_22.INIT_RAM_27 = 256'hEAAAFFFAAAAAAAAAAAAAAAAAAAAAAAA955555555555555400000000000000000;
defparam sp_inst_22.INIT_RAM_28 = 256'h555555540000000000000000000000000000000000000000400003FFFFFFFFFF;
defparam sp_inst_22.INIT_RAM_29 = 256'h000000000000000FFFFFFFFFFFFABFFFEAAAAAAAAAAAAAA9A56AAAAA95555555;
defparam sp_inst_22.INIT_RAM_2A = 256'hAAAAAAAAA9555AA6A55555655555555550000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2B = 256'h00000000000000000000000000000000000010007FFFFFFFFFFFFFFFFFFAAAAA;
defparam sp_inst_22.INIT_RAM_2C = 256'h00FFFFFAFFFFFFFFFFFEAAAAAAAAAAAAAAAA556AAAA556AAAAA5955555540000;
defparam sp_inst_22.INIT_RAM_2D = 256'hAAAAAAAAAAAAAA95555555400000000000000000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_2E = 256'h0000000000000000000005000002FFFFABFFFFFFFFFEFAAAAAAAAAAAAAAAAA95;
defparam sp_inst_22.INIT_RAM_2F = 256'hFFFFEAAAAAAAAAAAAAAAAAAA96AAAAAAAAAAAAAA555555554000000000000000;
defparam sp_inst_22.INIT_RAM_30 = 256'hA5555555554000000000000000000000000000000000000000040AFFFFBFFFFF;
defparam sp_inst_22.INIT_RAM_31 = 256'h010000000040002AABFFFFFFFFFAAFAAAAAAAAAAAAAAAAABEAAAAAAAAAAAAAAA;
defparam sp_inst_22.INIT_RAM_32 = 256'hAAAAAAAAFFEAAAAAAAAAAAAAAA9555555AA50000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_33 = 256'h0000000000000000000000000005000000050000BEAFFFFFFFFFFAAAAAAAAAAA;
defparam sp_inst_22.INIT_RAM_34 = 256'h03FFAEABFFFFFFFAAAAAAAAAAAAAAAAAABFFEAAAAAAAAAAAAAA9555555AAA500;
defparam sp_inst_22.INIT_RAM_35 = 256'hAAAAAAAAAAAAA555556AAA940000000000000000000000000000140000000000;
defparam sp_inst_22.INIT_RAM_36 = 256'h000000000000000000000000000FEAAAAFFFFFFFFEAAFFFEAAAAAAAAAAABFFEA;
defparam sp_inst_22.INIT_RAM_37 = 256'hFFFFABFFFAAAAAAAAAAAAFFFEAAAAAAAAAAA6A55555AAAAA5000000000000000;
defparam sp_inst_22.INIT_RAM_38 = 256'h5556AAAAAA4000000000000000000000000000000140000000002AAAAAABFFFF;
defparam sp_inst_22.INIT_RAM_39 = 256'h00050001000000AAAAAAABFFFFFFFFFFFFAAAAAAAAAAAAABFFEAAAAAAAAAA555;
defparam sp_inst_22.INIT_RAM_3A = 256'hAAAAAAAAAAFFEAAAAAAAA9555555AAAAAAA94000000000000000000000000000;
defparam sp_inst_22.INIT_RAM_3B = 256'h0000000000000000000000000000000000054002AAAAAAABFFFFFFFFFAFAAAAA;
defparam sp_inst_22.INIT_RAM_3C = 256'h0AAAAAAAAAFFFFFFFFFAAAAAAAAAAAAAAAAAAFEAAAAAA55555556AAAABFAA940;
defparam sp_inst_22.INIT_RAM_3D = 256'hEAAAAAA9555556AAAAAAAAA50000000000000000000000000000001040000140;
defparam sp_inst_22.INIT_RAM_3E = 256'h000000000000000001400000002AAAAAAAAAFFFFFFFFEAAAAAAAAAAAAAAAAABF;
defparam sp_inst_22.INIT_RAM_3F = 256'hFFFFFFAAAAAAAAAAAAAAAAAABEAAAAAAAAAA56AAABAAAAAA9400000000000000;

SP sp_inst_23 (
    .DO({sp_inst_23_dout_w[15:0],sp_inst_23_dout[15:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,lut_f_8}),
    .AD({ad[9:0],gw_gnd,gw_gnd,gw_vcc,gw_vcc}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[15:0]})
);

defparam sp_inst_23.READ_MODE = 1'b0;
defparam sp_inst_23.WRITE_MODE = 2'b00;
defparam sp_inst_23.BIT_WIDTH = 16;
defparam sp_inst_23.BLK_SEL = 3'b001;
defparam sp_inst_23.RESET_MODE = "SYNC";
defparam sp_inst_23.INIT_RAM_00 = 256'hACB0ACB0B4D0B4D0B4F1B511BD11BD11B511B4F1B511BD11BD32C552C572C573;
defparam sp_inst_23.INIT_RAM_01 = 256'h00000000000000000000000000000000ACD1ACD1ACF1ACD1ACB0A48FA46FAC8F;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[13]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce_w)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[11]),
  .CLK(clk),
  .CE(ce_w)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(spx9_inst_0_dout[0]),
  .I1(spx9_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(spx9_inst_2_dout[0]),
  .I1(spx9_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(spx9_inst_4_dout[0]),
  .I1(spx9_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(spx9_inst_6_dout[0]),
  .I1(spx9_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_2)
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_2)
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(dff_q_1)
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(sp_inst_15_dout[0]),
  .I1(sp_inst_23_dout[0]),
  .S0(dff_q_1)
);
MUX2 mux_inst_22 (
  .O(dout[0]),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(dff_q_0)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(spx9_inst_0_dout[1]),
  .I1(spx9_inst_1_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(spx9_inst_2_dout[1]),
  .I1(spx9_inst_3_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(spx9_inst_4_dout[1]),
  .I1(spx9_inst_5_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(spx9_inst_6_dout[1]),
  .I1(spx9_inst_7_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_2)
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(dff_q_2)
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_39),
  .I1(mux_o_40),
  .S0(dff_q_1)
);
MUX2 mux_inst_44 (
  .O(mux_o_44),
  .I0(sp_inst_15_dout[1]),
  .I1(sp_inst_23_dout[1]),
  .S0(dff_q_1)
);
MUX2 mux_inst_45 (
  .O(dout[1]),
  .I0(mux_o_43),
  .I1(mux_o_44),
  .S0(dff_q_0)
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(spx9_inst_0_dout[2]),
  .I1(spx9_inst_1_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(spx9_inst_2_dout[2]),
  .I1(spx9_inst_3_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(spx9_inst_4_dout[2]),
  .I1(spx9_inst_5_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(spx9_inst_6_dout[2]),
  .I1(spx9_inst_7_dout[2]),
  .S0(dff_q_3)
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(dff_q_2)
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(dff_q_2)
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(dff_q_1)
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(sp_inst_16_dout[2]),
  .I1(sp_inst_23_dout[2]),
  .S0(dff_q_1)
);
MUX2 mux_inst_68 (
  .O(dout[2]),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(dff_q_0)
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(spx9_inst_0_dout[3]),
  .I1(spx9_inst_1_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(spx9_inst_2_dout[3]),
  .I1(spx9_inst_3_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(spx9_inst_4_dout[3]),
  .I1(spx9_inst_5_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(spx9_inst_6_dout[3]),
  .I1(spx9_inst_7_dout[3]),
  .S0(dff_q_3)
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(dff_q_2)
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(dff_q_2)
);
MUX2 mux_inst_89 (
  .O(mux_o_89),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(dff_q_1)
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(sp_inst_16_dout[3]),
  .I1(sp_inst_23_dout[3]),
  .S0(dff_q_1)
);
MUX2 mux_inst_91 (
  .O(dout[3]),
  .I0(mux_o_89),
  .I1(mux_o_90),
  .S0(dff_q_0)
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(spx9_inst_0_dout[4]),
  .I1(spx9_inst_1_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_103 (
  .O(mux_o_103),
  .I0(spx9_inst_2_dout[4]),
  .I1(spx9_inst_3_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(spx9_inst_4_dout[4]),
  .I1(spx9_inst_5_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(spx9_inst_6_dout[4]),
  .I1(spx9_inst_7_dout[4]),
  .S0(dff_q_3)
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(mux_o_102),
  .I1(mux_o_103),
  .S0(dff_q_2)
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(mux_o_104),
  .I1(mux_o_105),
  .S0(dff_q_2)
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(dff_q_1)
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(sp_inst_17_dout[4]),
  .I1(sp_inst_23_dout[4]),
  .S0(dff_q_1)
);
MUX2 mux_inst_114 (
  .O(dout[4]),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(dff_q_0)
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(spx9_inst_0_dout[5]),
  .I1(spx9_inst_1_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(spx9_inst_2_dout[5]),
  .I1(spx9_inst_3_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(spx9_inst_4_dout[5]),
  .I1(spx9_inst_5_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(spx9_inst_6_dout[5]),
  .I1(spx9_inst_7_dout[5]),
  .S0(dff_q_3)
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_125),
  .I1(mux_o_126),
  .S0(dff_q_2)
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_127),
  .I1(mux_o_128),
  .S0(dff_q_2)
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(dff_q_1)
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(sp_inst_17_dout[5]),
  .I1(sp_inst_23_dout[5]),
  .S0(dff_q_1)
);
MUX2 mux_inst_137 (
  .O(dout[5]),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(dff_q_0)
);
MUX2 mux_inst_148 (
  .O(mux_o_148),
  .I0(spx9_inst_0_dout[6]),
  .I1(spx9_inst_1_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(spx9_inst_2_dout[6]),
  .I1(spx9_inst_3_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(spx9_inst_4_dout[6]),
  .I1(spx9_inst_5_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(spx9_inst_6_dout[6]),
  .I1(spx9_inst_7_dout[6]),
  .S0(dff_q_3)
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(mux_o_148),
  .I1(mux_o_149),
  .S0(dff_q_2)
);
MUX2 mux_inst_155 (
  .O(mux_o_155),
  .I0(mux_o_150),
  .I1(mux_o_151),
  .S0(dff_q_2)
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(mux_o_154),
  .I1(mux_o_155),
  .S0(dff_q_1)
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(sp_inst_18_dout[6]),
  .I1(sp_inst_23_dout[6]),
  .S0(dff_q_1)
);
MUX2 mux_inst_160 (
  .O(dout[6]),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(dff_q_0)
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(spx9_inst_0_dout[7]),
  .I1(spx9_inst_1_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(spx9_inst_2_dout[7]),
  .I1(spx9_inst_3_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(spx9_inst_4_dout[7]),
  .I1(spx9_inst_5_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(spx9_inst_6_dout[7]),
  .I1(spx9_inst_7_dout[7]),
  .S0(dff_q_3)
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(mux_o_171),
  .I1(mux_o_172),
  .S0(dff_q_2)
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(mux_o_173),
  .I1(mux_o_174),
  .S0(dff_q_2)
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_177),
  .I1(mux_o_178),
  .S0(dff_q_1)
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(sp_inst_18_dout[7]),
  .I1(sp_inst_23_dout[7]),
  .S0(dff_q_1)
);
MUX2 mux_inst_183 (
  .O(dout[7]),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(dff_q_0)
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(spx9_inst_0_dout[8]),
  .I1(spx9_inst_1_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(spx9_inst_2_dout[8]),
  .I1(spx9_inst_3_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(spx9_inst_4_dout[8]),
  .I1(spx9_inst_5_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(spx9_inst_6_dout[8]),
  .I1(spx9_inst_7_dout[8]),
  .S0(dff_q_3)
);
MUX2 mux_inst_200 (
  .O(mux_o_200),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(dff_q_2)
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(dff_q_2)
);
MUX2 mux_inst_204 (
  .O(mux_o_204),
  .I0(mux_o_200),
  .I1(mux_o_201),
  .S0(dff_q_1)
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(sp_inst_19_dout[8]),
  .I1(sp_inst_23_dout[8]),
  .S0(dff_q_1)
);
MUX2 mux_inst_206 (
  .O(dout[8]),
  .I0(mux_o_204),
  .I1(mux_o_205),
  .S0(dff_q_0)
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(sp_inst_19_dout[9]),
  .I1(sp_inst_23_dout[9]),
  .S0(dff_q_1)
);
MUX2 mux_inst_218 (
  .O(dout[9]),
  .I0(sp_inst_8_dout[9]),
  .I1(mux_o_217),
  .S0(dff_q_0)
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(sp_inst_20_dout[10]),
  .I1(sp_inst_23_dout[10]),
  .S0(dff_q_1)
);
MUX2 mux_inst_230 (
  .O(dout[10]),
  .I0(sp_inst_9_dout[10]),
  .I1(mux_o_229),
  .S0(dff_q_0)
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(sp_inst_20_dout[11]),
  .I1(sp_inst_23_dout[11]),
  .S0(dff_q_1)
);
MUX2 mux_inst_242 (
  .O(dout[11]),
  .I0(sp_inst_10_dout[11]),
  .I1(mux_o_241),
  .S0(dff_q_0)
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(sp_inst_21_dout[12]),
  .I1(sp_inst_23_dout[12]),
  .S0(dff_q_1)
);
MUX2 mux_inst_254 (
  .O(dout[12]),
  .I0(sp_inst_11_dout[12]),
  .I1(mux_o_253),
  .S0(dff_q_0)
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(sp_inst_21_dout[13]),
  .I1(sp_inst_23_dout[13]),
  .S0(dff_q_1)
);
MUX2 mux_inst_266 (
  .O(dout[13]),
  .I0(sp_inst_12_dout[13]),
  .I1(mux_o_265),
  .S0(dff_q_0)
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(sp_inst_22_dout[14]),
  .I1(sp_inst_23_dout[14]),
  .S0(dff_q_1)
);
MUX2 mux_inst_278 (
  .O(dout[14]),
  .I0(sp_inst_13_dout[14]),
  .I1(mux_o_277),
  .S0(dff_q_0)
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(sp_inst_22_dout[15]),
  .I1(sp_inst_23_dout[15]),
  .S0(dff_q_1)
);
MUX2 mux_inst_290 (
  .O(dout[15]),
  .I0(sp_inst_14_dout[15]),
  .I1(mux_o_289),
  .S0(dff_q_0)
);
endmodule //Gowin_SP
